`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UI4nZ9Ddw8Y+f646ARcxN5AsBu2bZ8W+cEBkb9DV4uXd0fg3SSDSnFfkYPqJFF9XOl0gi/rR09Ah
ie8pVu+4MA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PPVJb3AZQ+tHB1xjWfRQLT36feEDxfrOlr6rEmsPwLqo45vVHkw/jt9iOluxcp2SzCSDakdhgUsK
r88R7CQy+ffQYytnJ+uDS/onp+eGVl/FXoDZhPZeia+9Um197tJfCtxTr903H7kv5cuJk1nv34Ef
ktdNhCQj80m4S6jcB9g=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TSmC6xRt2CYGpDdpr5p6sp1lZ10hxMP7Yah6hn6Car4DqSQb0Mn7e4poVTZaIY/1V9VovuowETd1
eJetVlykUYVMKL4h/CV49ihzxzcwCSyAGg4o7CHaRpjrT1bqjpYQbCfD3Y1PNa52C/t155P42v0b
jF5JVfK+cmODby0R2T0gqc8K5S5ZAQWAbaiZhPndDCxftSg0O8c5z1txMsgiLDW31VR1BcpfGYZO
spOURUV+MLbX7R6AENAvKuz1iaUnIZoWGAMA9KJ5mosmeFYFA3WKBRwuJAiTKldVgcDhzaZmc+MI
aKH8LVWibbPg42G+tThoNGfBFvyh2P04HUjq3g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XywGaO5j8iNrlSTKoqD4L10CshA5/214cqHiUMk+kksPprztBB0k4HunjjRlJuadND26BuYitDGH
DkjErzgSAmcNYVYmdQ2T3+iwMxymh0iJhxihXUaPqF20bTmXh3jHqRsox9gtzxlmd+x6YkNvbc4g
eS6SAnDF/XbF22baePRiE8Js4V9CZbGbX+bVrri/2vzrU50jbBCjsUPv+BuRZUj7enx640mES0lx
kN2noLuihgMpb49kM3SxEgSX/A8I0f1xINyjAAlqrArl3v2LYdifKoRFH0tcRnP9wCFb0PFNndfR
JF7NboyWsTpeZ0iZCcNocVkXqs422rsmUHHA0w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aQGhZu5tQ9da8eMUB9Fm9xuw+YMoDIbos9IZH+SAB6mVeliAhtti1mKqdoCKuSgpXuCuUA53T52I
2Lub7WUHA8SBRPzVAyvqDvrjqEy8Uqgcaj5DeUiOBdWF7BF9qD3Riuy7C3FRw7qnqXURJCEvHuDq
Qws1RX1XWILoTr+vPVzSWNiqM7MyUyIjSHofjB4msb8hNzaqSjs95bcDXzEp5NTBqPeMOrwFxLoB
1aXHUvrYAMcT34ldlh5TOQUz6N/DleF3sJeRuBJSNuOo6LmUi0MJVZu1ZY+UXVZe8rERTDVnkjF1
ZLqqC3tXcFI20u7k+E9NDtdZpGqumwuNIVA9cw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P8GRuA18676HTrnJGqsWwI4RpPA4fp/b9bHdlLC5iuA/LXoj7evvLBkXSt7MSNrAnZaQGuzSpoc6
NAxs5g4c21x8vn1lHCZGZ3BnKu0SCNqKR0HUg98Rs4Ug7FiAIOIEFn0lplN/6bylgDqsZdfw178T
Ah9BWHjxxbJnc4RsNKM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pyppsGYHdq4VveATGiec98/blbAQ+Jq/t34XF5RT2yr/oVwbLEqs471n15PCkKz+r8B6jZk490ee
Jw8WJOpc/KR7o7QyeWhv7h1SHgD2STN7wY0u+3qNAZEWmrnKF0nhuXYs0iUfPDZ+86ClroeMoQzv
VHsluOdxTlB4Pvq78AWUXa22jRoS/SxJpVvT9ipT0ztFTs72lhGfluXscbWrZbaMCJu3UEXLw7eU
P20U2G0sI81Z72OA6XXrYpWzpQqY10fpvjSDCq7bxc7OZHwuN4Kbk9TYPrDwdRHwWNtzHDKk+Bwd
1XnmSSDWLwiAg5rmVBul4HCWHDNfo026e2ECxQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211344)
`protect data_block
mYX87PzaDZNdksorOiYwi/a+sOScPhR8s/uWDPp1RAZ57p/Oz4baEjIhUdi1NbWhb0wFYmzxqXDY
WLQC4WKahwnG18eC8hT+bJ39XmjcbDt0piRFtXNjfRaPFJlqaSe8OoO7vieY+5d0H+S94lg99Vst
FxQHciY+s+fDkFurJMqOom6xlIbeL0vGIbpbcDGgs1owIcXmfEbdY3YZhlnz4dj2/miLTAiEBhl8
7JQ7qIoAa2CO+opWPYCqCPa54LwDaL4Lzm27WhTGIHb4fwqjKygv7rmIFp7h6QiZ2H0yxqMuf6ju
e/G1bQcs9kUOmtECBNdSjpXZOfSuPtUp+Yu4yiEfIRRo6vyAqPiK8FwQTb/4lnjVKgorQmtHQqZ4
0j64YodeabFV7t8DEm0ogpoFYZYjE40e0kYwcgLt1iTHE0e4BXOHDsWKq1aNwymKoknWf0jJssJ+
5JIrXyTRsZLbWwex9jnOmWVoqrcoO227msXs0EhEtXA+YXgOdt+z+Ou8x5XYihboJbBHJ7RKHGig
H/OSbkquyTzJhe4JKv73BsM+3GuBndWOuTA/4koSXoK0G9X0PmIE9m1AKowodOFWq8EEFBQ/cUod
mltA5cLjrCX47WelX+tFOT5RT7G8EZUeOIW0lNrB6FCoPouNioS5MxiH8N+VRh3Z/jr0hpOh0KqP
DjmqYZk3IH0jTUxgVB0sTTjtViAkiB+2fCMpOVAl7AQOlfJQH3RqeHhxYF7P3W8CnFjpn07kMFYV
bf0/eDOHXV6LYJ9oFxgUFukIqjpaomyyfwJBycgp+gAbKIGEBCSzhGiS9CwJ7yRlYFIt0z2arOGC
PKynosc3Vg0IcK+P5bawZXcd3t8zUuZ91i+x8us4QocAYAftHsiojUVaRd1tSIIIC5tSVAz1MoIM
DJidmJYofOfnfVDH9xZBNNmAHlftHeT9aJ8U4buh3xN6T/k6H6kMJa3szxrOF19E6wr6Sn+noN7C
hQW3p0ppevGYvB/FAj6ALT7JBMkBudKh10h7EEwLWZ5AfiTtKtGGhRivAcCoW9mEGLnygVoaaVkI
JkxLNbsDzH8TFcgaPAsTQetCdxj7jJuFQJYYhAyEyYLrfTTKLuixvgqDbrNqs32Q0M3ZTK0akbjB
sFduBZ44YzENfd1ClXfdRW1LNW8z8J/vryKdxIp9yZggXqL0NiUQOaoccN+Y5XEtXJzDACHg4vU3
EiWr1IfbpEIF0xs0eEUpHBlYhJ9Fi7yqnLMKNDIroDZskOKJHIOJYwks4bOuE60aTEdH7ZaRPEdk
ClZt4oKh9zpDKSRLyxw9B3cn8hBmf0Wrtu/IvqH0wsNoz5NVT/lF57tEKXrvvLUjArtA8hv7jNRk
AZguwtQr9tkK3jxchPrq2G1wZKSPSNL3UQUsT+v8Z6k0vPyyTFUpqu2Elm7tDulv3lHa0LXTyIm2
7VV+uh0/m7KvSACzB7PRxspq8VQ+etitteyvNcp2wDOGAfvwet1goS6a51G8FzO61jNKlBaM4gV0
OGtySJRr5FLE1JQua+Hcs/iGvZc7MyXDW9ZYdpGPV86ZoduTZLF+OSCT4kzgRhR41Pu9iKgm537W
BnhL8EIFl6c59VM4xyqhxCk5RXYpT9MYVGF3H97c/uR9oDLNvU5t4dSzW3n/zNhYwdUzaOI34414
RhRBIp5CsJgPmT2e0h59Oc/sr4cRnkZWsjK4cbBo3/EzgjpRGPaB0dm1TMKXoMg0ukqnWIgDJj1E
nWoyrC4IaB/z5HLplL/cLk/b7xkLuupcsOMvCHlpRo6+TfSxVQSW9fMJ8B5MaEC4yArSIEA6v41H
fxpmTToctuvogUnT8n56ZsM4KlXl9wEoRiaGMo1ad8z0QwFJQJ/Y0Z+NaPv7P4Mtb3diSTn4v9cV
IQFvKuW09JZla3cdxouZidjM3EeATUqAfLPaWNSgJlI7CnDm1o5wnRhM62KV8JDuWwlOfyX0Q6ZW
qZ2TLp8QmwWTDhH6H9+Y9j0gyX+FMRiarOANtxCqbS3aBHgGiy1dB955F5o/pBAP2jMSaACpD/fx
9W7Xg26XaGEOTDL5fYBNcE7Uvx7XWOzeKwfFKQY2vC9bQZVe4B7RTnBTavXKpjW+pcs2QBEyHIys
5im56eX3n3Ul2/zwisi6a+AXKJHfVJ99+2WCA9vBNoYR9CeRKKRGvou7dmP+brBwo3bpcMq5Q+H8
e7qG6J4m02GBYpoJ+s5fASX8DHm9obh63vmxQnpX8aMczVz/cRcIg0WPeRR8h9wuUlALE5Fq36ok
rWMVt8WnXFrsz9vhYJwKvNBVIJet+fN+dBSlerfQtfzzGGe3qAWOyznPjpjMmYyjja2+eXjXoQ36
/4LsUNmjY7sZ1IvuAKyeZZyFBESL3FtbN/ZV0sCniU37ks0ymv6TISXCQX34coTMUNownX6bbbim
iAAfnsFRb740fICmGgQY8AIE/SJTKf2lDuBJdaw2zX4M9t8Ynym9y/ZKSw580ffy+03dYVYgPtq/
bdihDIKJdx36JaSN5qW5YgKOqDWpbpTnQ1iBj8mE8adVf1SMXub95jvjYMM7mGYX5KtdusKHuqr/
8uJ3Q6uFjRuDZcblSsEUrSO0RtOBDwWNcHpngQ9Q/jv/3FXBk96eTS6d2OfhzTkYjzPlFIgoxOb8
MEr/9Uf4tIY+ogM+ndGAR2ZD7q8LspGJDqS0Zve2kO0wga/Xqm8n3bSAeaJar3M054qjSBZNLPHO
FtTS/Y2zjBnNjr2W7U6RCTKw0wh46CJcNL9qeM1tnh+mYS2gHx8NRV5iAvvJbO7gGzsl7ueQu+bS
w2TtpUdCNO0AJZBfk99knkClKnPmPlENgSQMhFT67iYEeCjzMWMunpmdQnBh3E3gdofO/gZ84mEN
LcEvXEu/p19IxWywui/L90HWPaI2tjjo/qDAM1zwrEvE22P6O+58YJEfrB5xLxyAyOERI+rjxIz1
YUXi9Lqz67+cNXDt4OvNfR3miLXGUrI8BrtAQeTiGwNrKjCP3w8G+hvfPuC4nfXPC3/r1ER/57Bu
RAR+lAXMcN/9BR/H93CfiHZhem6NahQ+Z6JxqAkEDbEaGO0qiVXRPOhyhirPeuNNJCoH8zbYjZg3
oBc9x3Pd4DCD3xjguXGIltNypTCgB3wYZEQ2jaYbywnX2aekRbssWfkeAFj+9hpmNH/tB9VcD6wD
JUakBbvd9VSALgTuYa7sN13r7ZQjPWJIQ8dohigy5pYl3K/gWRliE+QT0L396QlJld1QjeR7hG4x
xYH7rcHvj/qBHmcqCL2vqhekZb/Q1z4KvEUizUWoltXuFv73WRW3bpksiQPB9z/j3cZ1bkjss0z3
h8dHhcFGzgIC5+/e7M6FIaQr3Lh17rDQoa8KHUabdYD20DOu8eca34G2kkcBlgydt/RufUdCWIGD
iT+z8WiE/bZ5VeTAGxpLtQcbsnPIgAVEmSeDEJpfAlv9iXjvKtipINyh67IGDzYgKWNZfCHNaK+O
kd+jbNL/Vn9KIOEyul6GhZmtyVqErx8sq/blDPr3hAAh5zqFiT/6M7YeFn/AIRwlERvCmO9nOC7D
9Aebv1lYCtY62KwSkQlP1qEVaXKSRhHHh/M0MeUW3hE1pKYGdnhrXTr4AeeVXvjAs/gzCVrsntI7
JViFqe7C2wskVXVZadYKBossqbuYkMzedwnSH7rfxpnOC6izZzpGL1OHnyke7cATP7rQ9kfeW4Mw
smBMI03ikL62uo+Rqru5cyS5/8uI43ydHCbYa9noqt1L1SrEH/dVpSDPrHhblxUkk+wZgo6/Eb7h
NfSsVOgRF9+Hkz8z3ZYqyD/pEBsdcoGyrO3frhwHEaBlbe1JLzWHABBA1EfAWpw3WcMhO74kbHfj
FHthn8UVOLliwP3Qj10ZfUxrBI4r5bhSpMtyiZCGjzkS5Ae49V6qMuknge0PrrBZ7Sdlec1JcSqp
NzbJX9HdTgOMBEcT7HVK31f/xRr1bVyt2pDH9MdshPkFW/lImA7qbpqxQDSCFgFOZMV/7MiYKIDC
oSPGuaY3rGTqaLkz7O0qKx7Kv3kQonx2G51S5PFUOtsQLuoVhOiBPoE3ZRGmJYcwzCiYnBpgjUer
fQhXUo9dsN94vVVOL6kriXwQkffKQvEDa9pPQtfGPtZx7pnfJrjWSf3D7omc06fFZRDU4/5rm4ab
RUQiaRQZwF+Smyj7b91a73MBJlkWC2owQSrF86zUyycpDvE4ebGHjSgQYNbkI4ycZ4prVwcAExzL
hIIoLuUiCgRdrBWHOT2KiWNGU5YhiHn+zzlObCGMsW1HCaheX9w1YMC0JMWR0TOQVrLbwpfCuRzj
MJ1sV4gphcHHlU13v9kx9enr3N4ZZauOY4hqE4neP2/FT2jV/lnCovDzQ+sh7q23BMeWQqsZOFpX
f2QaWYZOkAcGLPc8iLw2BiJmJqre8+b/7CzLBRYlGtbP8Af7W+BXEWNQxDRpcsYm8xPOPQSdZrAq
VDddb8EzFwUci7uPsT7iKbV1FZAWlIWcVfE8tIVO2bQLcxlkESIssmwU/6kZxhxA5BPnaFWe/Bn2
o0DYRgQzZp/89LFuSOl+047byMu0DO/GGfATvbwsaF+IREe9NYdgKX3NDhEjs/mgq25NCsbi2bvF
yVLJ21KbcUtdGjVzvyOZB4nsHLN3f+M9x3nJXqDnirxD1vOQXA3Zl7sxyzL1zAfEkZ1dHLbhjN5e
+Ab3agaO65D5BDC5m/hUVWGpdCI4ps1J29NoE8rGPaUv0KCGd71LtuKci4elRh59VpgfwxriHlnZ
JCU3jJkD2Mh3IKVSLIVX1SB2chIscdK6XgAT4vekiZyVAl03Q0nX3M2VKkYhhesGGiG+o/Yl8XvL
pQeo3GPw/YHjmwUVl3Lfn8jokz/GETplsOEHzZvOMnvZysffArlyvKPvljefnJoZNsOBhfS5jYGP
hQaa/xSQ1lVuMrZLuVIOhMqTrYjNCtQ8sIipTgw6y5BJctNJeTsgisOXQRytOMCRCvHGBZbW3PVq
n37kzm3kEgvO1If5OEocuXJ0JngxITWNWID9N+hPQQiZSp+vKQSySYfN5kNH/Nl2i2CbyWNS12l5
UUlCKKDbZvp2FJ2oV9n1HCiQAmj2ZIpRann90nMg1s4nCecCJh6KoEfwGv4udzQ7M4icbB77Uri4
ZiqGdTGase7gz2pqSMzjwOWmlr+Go7Si39p/zW/rz0/nfmWJ0WsvQSp3ms5C7mjIoiFvwGibTsqU
6q+lhTS4f+S5Tf86MwZRFtoKNTE4OCq8NJ+7xKgTmEe3XnBjGIPH6hEADtvtUPZGpcQosyLxX33c
XowNGFIx31VBYKW42VTTYXQPqjAknwKyJftoIYw1L8t2aZfga9t0xHC1BIbVxdTGrxblT5sZVXYO
MOGWbu6ZoMmUydn6NI4wAo+/m8xfdlNn9lvojrRs/v000gfavAAmUkHwPYMwEyS8JcYW0qh4jCdI
RArz0hbRWa7YvfLrem6UKyR+Pg1HRpCpFj63hoaZRhevN6twz6GvheSl6ZZD0j5HReI4BJ72iibS
jR2mY0NzCZebXmBOTcTvQQkCRz3/5f1suDOu2gxY1Fg+nEtroza2IbPpAvyMbgTRXiRffBLzpKvH
W817Gyuy2NIFmVZxdLdcWw+n1jDru67SP+CSggD2RVAz+k+ijgKGLQcGL4tmFMLsYKN6NuB73Y+F
fzlJ22zXvvyLDEV2Lb2Ch1AnrMs8zly7iWS7dR35c1IQjywhV5n+fWtqfHuxebT7PJBTmKUbkPTr
D3dYxyqcbr7T+1POLUVkYQmq7sR9Vf8yPi40KDttwgbhD0qDI7Rj2+itpohbHCYdXHGErEKTDb44
hZ/mypeXHEoTWfr4/g1dOJSqKvog1lcU7PUeWKEHC6VSyaGnlYq8IWaIAzSMiTcV2JlfDcW9ipJo
oGcxGTceSQCeAhnlvaccPOL2Mcu6SX4U1vtIkjrWsLYHkPmIwFpW/ek0M1MINjVrW0nOLsuJFEdq
CAFWnKiZHQobhxNZDL1oQ/WZQMMsUafJ3B8rAoBnw33tHzgVwLpskVtiUIm6q6ZgOfLKvjfhGc6o
fbLSkIhPJf8tDah1mGhdZQadhEdoEW9PdH6Oda1up8OKqLTjW35FkmA1hzl5rtiKNi3aGnNR8btz
VJJMPqsyo6is9cMJl0usAXovxNZqSa4U9okXMo4rJflLe4t9T+PBZsICR0tw1Ep0g7nRfCg8hmSc
BbYxqfUBtbOcqyAEuVP+NTmJowzXPOqkrU3MsY9BhnKhh+Gi7mrRvBtRZ2HU0G41CfwWwMKTNOYr
L19jnHFxZrODYTjjYeesyzMFzf7nMwjrIo3SIupuYkUG9sVLyEa8QCpMp1LL5sQGzNJqHKuD0dGw
9RnwHqXKdPAkAbBelSyEZ+eZprdJWevzdYyWB6j8voNTR3WlycxsZlrw3I8YhwRQVX/T4GhMmSFB
2WcUJ9uFUUKn+J3QJ3oH04uUgR7FEQGk7584rH6blVRwIeWUQAx+leP4LBMOhz5rzESr84lLTzBd
FIh34rltIhESsNaF4VpMHfC+VWeeqXGo9iftm2hYktGF7zpMbXXHWhgLp+5IfZ8YbqnSOWTfdoFQ
GOjpQVy53QQrt+XnsrGhCj5pM3eLfJrZLmNRC+TFPVMoKFQDLfu20GkRn3NvX4LP0kC5PsWGNVws
j5ysFSS5yBgxYLI8+CCaSxWMTggBJxCo5ZEWjZVzGZiiHLVMLdyI4qIEpQNsD7s8mxTS1OzdTW7Z
qs3JBP1Tjo8AmHrson33xPOyr1kMIw/EfsuZ/49Zhk+/vSdz7ac/2mPoNwaai6kNi0ByREqnA5U1
4pVQxTSIm60Cw7H+Xi+wclhn9kDr0GcAuRuwfx4IHnFFTnlru9quLY5iWeIaEzldifTaHyPpB3pu
xRSgpdYvIopEMzMD1y8Hglfx8x3zNgErbK1UNk49wwmzS83L2/CxJMj0CUfrHfqGd3GQAxkRgLCf
KcyiXLb1gUyi6XnFOVkIecFH3lgUnMmUtCwS8raB5yK5IsysJOaK/wyllrMqHiK3XGrjbQRQhPHa
8x5BkoCZBUec8EQtf4A7iDczKMfvFtLXszMpW0NaS4ZuWFjlUVntvC/irm+l/JrBNuM0G0lyOheT
bD7tlECGuU1DqITAPZOm7kxbe8uw4/09daRONOUH5vua5JSzNIc+gjMrCKhbaQdb0kz0HcPB3t3E
tdgJwGHkQF3LzeWIMtmsQPT+LqDwM4CJCUPkrPiLLbeg9BdlCPfyKb72lPsaG83332lh2DxPb9Lx
He4CPqLDkX1cqusAYHV5L5v9RdZC19Wc03/nziflTeKNJ5DJAouXDUKIyHX3xB6IZRh9YRS9WKD0
OyzAIkMpZ1npXYGo2CfGjl0c5WSqoxaku6VC2PF2E/tbfVq2sJ7UGzxm6IThyjPzxp7jvJIMiCRY
j12G+FU/DTDf7ycEYeG9IEzu5jZH4CiYliafzsSHSsDsdVWBoFCXm1gHeoo8z1nMHYmPr9bfQhiv
9r/rumM8fEKwfCWuLj/8sPTIh0Kg9govqks2M3Oc64KmmucdPm8QK7xvBSDWqD55BQbU5/Kd86Yw
Z2kiZcTvIypcSHyY/VOFFvUY1BTmWfKrGOkyyQeqec3FzH5kLdOUYp8IQXLKmDWahTKnVKoWCi9J
1ba8LjsM9W8q8Xtit3hn6IqADvvmjL/3MGPs+u13zZIkuSVgH1MhwHUZ1wWNvNnc94jDIy1V9Uub
NAQBuKRrUW+RIGbXak9VJdHvgjCej2PJnO8plXfSSWo47wHhBZ0BNCJaXRVJNB8RjrDhb2M3q1tZ
PQvDAKLsEbly6mgoUhzCGIfAjusEBBQIfWyBk+3Is46xLfBb43pWIIVYKHV9BOGAJKn77CdoWaIC
3d2HC5fBRmwaZhzH+z411SFg9NiBOTbonYZTNQ5dHD717zHigVQFbKyd9vNSTcvRBC0muqV4C+WT
rYdo5o/doUTi5vNBcVJ+IfWuQ7Wv2g0fJ8J3ttcsBlMMLXzmhExUM8mWUNGW08GOudm8nMzCQIkJ
44a71LT6ONITLCf6NnayMIjg4zJuoSE3Ih4meyKEN9biUDisLJ3gY3d5G0iYwq69zeiVcuZ+umqM
9b9lb233zVrTh44PpZ15e6MDG/3MR8mI4Xne7x3BMypHBLTbXgi9AQHuEoTBU89oGT9M/M3U8wgH
TigVFi3zdyoTJbCVIMk3RdAcnS0SoYM+vFPAsv3j8REvp7xK9VGrCVKABwT1mtkcpr/Sw/nMoYqP
+yD0Chn2ouamWhBnwRpLYKlt1E535c0wBsQ/3i6eUo00rD2FxBa4Rgrk2ubzkSWVMWWckmNfn9wA
Y3ZmDP+juNvozBfZDTIUNvEix6+8syVU745t/gsPZT2oGGPt/VfdxjwngEyUhTty59asHu4pJxv1
k170rNi62/FLAqCHfLGea7QC0QJh04BM7joOXZIjSl1yz3AWRtglq4Jf57+O9qZPFEBJYSx9SwDr
ya0xb4rR9uGnj2CwAJVkHe10RB9DazwI/B4WRUXqbrR3qjhcxddHrqxuZuhNSJvYV84HpEglMnOi
62fsdO6jRlooRQD0DV8Kn7Ir4EL+0LVPE2QFYfDMhWREbKvrxf5fyEHM4ot9m+TvV2ZsiXr+SAP2
HVbysKU4ogI90iG8v2xoFAQ/DBZtusa8DbixvhkgrU5/BrNryUHeuHCLYSqEubpxujlAE40eWdPR
o0dPAseeECeMUTFQ+VLznA40DVfY+vdEp9PgH6mM/uL1M9wIWykpX81/yOEEw9Z3HPnqBUoCwxGZ
i3m/JVBEYpM9qdWJvmD04g6Os7oXP6Yx0byXx92s7/ZkAUVD9cbSOtL59E6y7FvPrOn6iN/j1VrX
krFLxZ8esMEfkRvl60Wmu/PXFP6SsVkvYGaVZRiGLmeTrhIbTxttFjaKNLwaiuGoG54AHV6E6h/D
njmpS+tYBUK6YXkquleeGfyfe0sXe484z8xRBt/hYuHSOdHUPCF6UuJNDc1zuuAkJtsxQYx8WmzZ
x0BGMKZhwBu+a7ZRiQGuEPtWORMsHTQxHNQaRQEKXbehos+16lCTIQBcm5qpTaIm8qBJ4r9XNt6h
+JsxkBWEhSHwaRJw/rUwIn1pIle0isB69Ow2nWJ+QQzsns7eZNZ+Lp4Wq+HZyqCweTT2MXknQ7tz
oL5JqXHYkSfpz/f0nZhLz4mEBEJ2N/3riIqhlQ2OZGWzKGv6zlxiyHkk4KjHChza4psAoNuCIFK7
RiPVJ36CUfRhQBLxNs3IP4RsO8Jwy6FQHv7ZMXvDqRQmCpLDDrGPQVGuI4xrAMw37gHltd5zGqM9
+o8Iol3Qw0EwjMtFHjVIbL+LFQuTlgHj/E04RO20D51sFk2930Bv54PMJTYSW8WUK2hC2mVaRkTM
URJ+miU5b1dgPcHA9v3p62tvZ7WP2/QOIReLXele6Cuw6AhnQEYRwxzuuJWn0UBA8JguQQy932lX
g34RxGr35TGUzU94fOCuabgKXzltiKzNvnKRFAA8lMFyqSKtLkEmYXS1kPmTi1I/Rp0K9Cz3YsZa
LOiLzabkHzw5V5z3zDnhDQ9eVzbPgfHvj3TfKCVfatKYTop6plFUn1nxEMxHiULjrORec5J8LNDh
6JSoE7GPTcqm3bAoPonT4ofZ+rbOFsITPMqAfKu2KTwXerN7rELDbjNH9ceedzxFZUWPrbCLMzDU
fHhlHQ4oc5M6md+3lwCCTRZTCyKff30c4+kjNeLOeLoecbwXLiShaR2rYXKHwkkwEk0fN/lp15u5
peZQhGG/QuSHBZ6FxxJ0bXODlW0glMCyL13hnDklnOEpdm9ebuYSBCPe7XXJNOXw6rt68kgOU8cR
BPQwP8PUjIeWrM4Nb3kmZlf0x/mnuATYrzvMqKUGE8iENaj1uTYK+PwAVP7/v/Ji0HC5B9Q731rY
2Tn0daSvG6JtCxML/eVl47AdSkCfpYxAjAW68PFXN3d7xTUl1TX9L9kSApOLdqZq0Il0HtsSYbB8
l6rXWZt5mG/yi+5GHYxYuqrhYE3pxdGlX95/vwDQDMNTGYJ+TmmWQ4LNnIRp/0ypJmU171UsXYqZ
w1todGkO/1/TzHuHt8PwqHr/m7sS41RD/tnVjc45OrOx3O9e7ld9fhiwzoFsPlnz2gJgLIMPX4Lo
Of37SYMs0H/uGg+qrO35S/2txIKDsunmkf6XKkY25FxwholrRw/NS1rsV//N3b5uzhv20EJDkPHd
pIE7Q4ynKV1WVF1KiEsxPt+y9WwMjWhsHFz0Z5R/tafBGVKddX34kpWA9WAc5ShX3JBGUghIkquH
UWmEN5yaMsQ03dv6ozBEGyZHysOzLvzSJWTKbrlpdPrXRaurD0ch2SLH6aYiA+k//5A+KdeV8yol
RCjjVGIXaG47GTu5bg5iLcYK7rwhyRDGWegOkg/rEEUxPd0uG0nYI4+5XUuaSi+ozHvj63FuDCW0
VCKuwn+0UjjC78NRx7dNIi7izaZlv/7AyLwnkUZUAqlJ7pnne4E00Rs0zWe0Z7J93NgbP+9WMRMe
NGe1ROmgLuvEO+EdCuoecTQusAhNZVbtBlWyFFR47VnzCDphZQT/l1StynAe/GIDfvAWtN6Kn2km
kh1QWplQI/pRtZfeWUaRbZi3+37OAFhF9TFyvCcltj2kx85QNZDMtbKest+tGQ9CajulDUgt0bEU
b/wmtNPZNWjMpINp4dh3fpaYgfAL0eyTeY8AJ+K22K37D+5YH+5RKPnjI96/FDDAqKPx32945686
Nbg7ER/d/2mREdi0Sh+3iHhZA1Ix84YzYMMN0aJoOACEDU7c7G7eIdy6j3kiXavuosA+cPLvKEsJ
EgJzq7r3zt6DK7zOjnnGKmfYwWoB++aThV+yuh2XIPvsXuCnjUb5F/jipHWz3UG+AnqG5sCpwEU9
35tPXE8a8cvlf2PYxLCbNElmo729lGlMwEL+vEIWbpTrRjdcqm9cXfV5ImkefYxd+GJMGvBuSr/r
M+e71KiTTbP4Wg2fT0LIrbGNwkQa7QjbCKgxNj+xx9LYEwSN0l22W8G7lAs+GILsTxuaB/SOvI9c
v8x/J26gjgzTWs/jtbcY5DIDAqJ3x93w02UU7Mxq/Kn7C3P3LSCyyCzkSCMMU7pFaw0JooZPw4z1
fs4vnaPxydKbM45VtD1odbgGEOkibCe6G7j57n0r5Bphqh5era7iiuDZ1jg129iFP4K3bRve0XXi
2Ie9YNEweXZ80VGjJU+JJfnb9dw72WMl+LbtpAJ5iL7P5Lf/OpDB3/dpnrb5gz8a9BIXO/12dpkF
VxVIy/rVfU2LlW4Pft6t9j6u6R2DI2r+tZ82gZZh/i4xZh+4ZyOG6egjXy9OeV6RVbnpOVwhuOve
hZQ4XWs1GfIRYX6e2XBylEYGC8MqXnofxIoa5eGr6ZDxQ8BSFzHqYpoI+CaIz0Bs53ZoLwGH5IpK
KXj4LuTw+PNkj0MucxiAC8m2icHGPMIwBIfWgGCyfS/6z4FgG4hga1cwrggZ/wreAy7KhF91Aadr
qf1zSU2TWHybTGPlEX7dQONZ3huD3H07smXIzComQo0AVF0xlDUtGZbjOaevEzKq8BwhQtqWHEyp
BkD2OBaEbrkphuKe42zQ8NZ6db+mJNodk8nD8GD+8OnQcT09rGtP/uQojozfu6DKcEkdg8Z6gdv9
cHwfjtZOK9qIWJnLPLSmn5aw8tKJHVPDzMNvfBdiF5bQiiqankAR9GKBx9lZKU2JevUHzWKexozC
/tvFkn4IExV+qeSGIosTD/Ga9lkk6wA81FbCd6ObS+LT3GUpZXM6P9ltgFAbYvK6ClvjgLncVVMx
pxNN4YkMa5ka0oe/I21/U+EUoEy18Uq3OyFXvDoQASjIPLoSATkqgus9yt8DLHKzeQMRLGhEKr9B
Oc6ah2xAU4OUuroU4AaTATjaDa1WQyPGqBuKD3kOnAx4g4xffDCl96zWeq7RTDq732iljU4g8JyN
Mf8hnqjl+s6ewTeG34NvMF1r38EwIspqnv8Wv8K5OJU9QNAZ/DX0RnPhEL06KwqEe2kW1zbfsQ7U
E0dNMrkj4pwfm8OJwknuy1Z6TUxt72ABP/lrdCVc8vfOG4q9V0R6yYYLyEfVhQ09n6rVY2HoSlir
bpHhgD39+7L4usg+aHp+m3dNuWE1Bksz1njiUOiiS2c3N+QW4GODh9hlk1q7Y5Usdb1zWzuDWJkE
IvQ4edOZ32Qmg6BVAPhwozguy82/eF6sLIaINW8UNUE1EOYRXsQ56bV/iLWAViyhbw9THOIh9ZlL
oZqRByMrROTeOLv7YQO0ZD4Y5wBKQMjy/xw3GnBoFr0L4KRAqoXHQ7VN9FH4Aj7+Aa3z2uen0L7I
OHcAyx0x6ypE1MEWLc5AHIq4PNIYFT+uLUIf8ekR82szS1gNgRhdxQX7vkGVTnpYWiZHZ7IKgZtD
wq6Sgg1NpmvuPtT8vD0sYYsxgVbVRFom3xMbgSKG3CCe7MGXj3INZTZkadcWeBIkG7fXJOIqMI9O
P4OjF6plzZFKtD1dPcqUqCjFjadVfVZO5iT11u0qqTQFsuNG+qCqOPN15+jFe+3mHGKGHZwnrqIZ
uZ0t8uhyjRavnBZAa0a6crqhW1ABtKD1ccOUhtAq28/czSow5XP3GUM65Hi7Vmo4XAGjrJdSL7qG
Qozjs7n3glUAGaVhngL0rWP/i/hatCO9zfqhYVQg3u/iuHRV8eTj5OByxv91SYjYYPOQawNsnZ+v
gvqIdk3cSRBPeGjcEL1HJOXqqp1LD7MIUX1xHpjuBNYoOOOBCKKpxSzQDDKMMTbzTvRvoYW+57ma
RmCfiz9p1K2DCuftIpsfG6t47ffuLydFAnZReDUMMLmXWb9bBnpn10+0u1Qku7XgXY8og6DaQggs
oqeUdjiLldAwx4wWXH9UeUxM51d8O3pGkVDZEuSdtoZ6RkV1fWjfDCvWJMC2Wj0BtNNsCerOVjY1
6A9Hq+a7I8CpA2hTapovDpsieYYm9snnpGKPH7KioEyEISkqcnHNDctxlzKxwtrcmpeq79vhfa4i
wbFstl6zMKpwfV3YEkkanjipf4QxEp0ujuRP1uY3fCdmrG2lyhabpGa5hyEpGdChuMOTx+NnbPU6
sPnQmlrCaeeC77cO6Za/Dk1VPaHAY0XJhB2+aFQpsF2Q3aWMdxM4HKC538o/XZ7N8mymmYZ5TkPt
jrJdKNP3iNVfFt6cRgaza1eofJ3VaWIXIApFxFNwssazotrk9HRczsr036hcnCgpskRiAA+OOO+H
9+5DN5f2JU9TMFpJPW/qUERP89KBHMEw4UZFVTU1jPgrq2NPETfpKV4HAy73LEFRXBjOxTqlWIHN
1CVbaDv1Ez2yhhhqS5zrES7OPFdqD/Ic8glSGfII6HDjzL1fpO0v8KI2S6eyG17OxcoAo+y2rBX7
62wqhF6+CEFYV/yqfGrYlPQWn9tSd9TBHbEK+/HOmaOSPRoKHA72ZTnuPi+eznva1haPubImllit
ExLodMMCIaOhav2JomK30cxHimPVpQ/gUXCTLl63CA0WFX0SZPUsEi5GCC1Ej0WKGtvp+z6bsqhR
LYeor30q69tY35ZD/zgZ4eFPVJ+Lnvgzs+KRKsLUtnABFUCk6+ulkLX8wmkw+R/tUsfxAuyRw+sy
qC0iZ7opZHA/uTNJTFFC6Sa3kzyam5d5UZbzo6JUF3iC5GbdcuUANQ81v3lcjO1cqn2bVwOQEaJy
YuHn1KtlHQA8ytwbqjfCbqAEq/FqUZyAAsguhG0PY8PGjz9dIqs8rxFpr+HUHezrbze2iJX8yVlb
oBDVnsa6LuGCRg4YeueyxIVgSSAkZ5xc1tXki996opA801G0Vy6kh4jkZXtU63U3TkFJYj+HoyYw
PvwvBtm2PW7pdGWUUvmjmOW/9RZyRis9MF/6HuoeIUvTzRsZa3VbYKdmhQp4wAl7aYPxpopjIel5
ko9Dfhvz9PX+HP87mMzkvy3v83oouwD81NHoTit5haONbQ7PS5C9e5p682CVRT9qomvX3xbN0FF+
XcxmLq1fI2CiO++LxDxyklN0ZmuXAFWWV6MY7Hm4l8WLk9h6pxmZiDpOsyJduL6IVjLdiG3hZH+j
fLoT4nwySgsvmtSPswWiZMAGZennR5no35CD63GZ8Y/43CvkD9dXNsECiW3j6pgP+mXRUdBM2MtN
mrnjIi9SaPi2Vcmj39+iYjRZ18uuM9n+onaT631m4ShvE4Ks6acvq1VhclByoM2DLnZhej2K1kd9
cS8MD477WimDcdf4eHkqR+XEsm51+SOLYSMJYttxcqRVA9PIv6+rpqB9KJFuycrjluf7SBq+iBSc
qMbxBmiFYxFQ5ynPFYfVdr6t1ZfaKrffQ5xL2zxve8oIxKRuWoy/Y0pnvwWawB5P2KrDOqc+p88P
bB1I1wBPHQMtwzxP0e6J/jGPodmZqTS4Fw2JrGilZV5j7LKFcRyfPMVFjoj/YmxFyyArasLwZuMh
runOa8bKCd7TBTEfKxX4XFv/QIB1oh0mp28auM8YHq1JwxOej7LL/UgP7ikWZRECjhY5P1Q1LnjG
nguuENrL1cMbAcE+Br+PVyf1nE9DN583p/wdjBBpLUR93VmzFJxIwq5OqgE9c2qftkK1Nq/zNq1q
TwielhD4cvtySZ7apbll1/3Zlf3iwi3MoTaCPW3jGkpwg+jf+UwLabLZbhtXrvaCje0uQOX86+UE
FEnB0Wcp+kr0J5zBuW2Nr8yGJ5allLIhi2D31lJnage48zRrCw9Dcuogp3pelMVQnqtCrmwrXZPu
ScMDbxN6/8S2B1Lv5EV3WFkN0i13cqOWwkr/tb9WD52HaJzo4ck32jC8Loe3qEPHMp+y2FQnDXEG
0R8vlkJnYY39hQyEMk58m5UE8pv7ZC9oNok4gnDZ6FleAYs9az5dq/XOIAuBr/yYSlpL5Z8mtJfO
Bke6+BLWWtTTvdXrKbIJhqiD5YvvAdCv6heO45xvWmsJeqOv+ReJ5XPevkv77AL5UCJTKeaWpwbh
TR1kkOlId8XV0PBZ+FmDDUOZYKZKPHTO9cVPGseUhUqCPYFk1KJbHOVsnN+cKxTy50yFYch/FhSh
IJoYPHLzjVxAcjTuAZNjrkVH8noWZzdkkx4UiNUV8lEPKOqKubUQTBhf4hvWSaaK+B3TP2MemrVG
weq4Zpj7BIvFTjDiiwQY/Yf8Syv+YjYlfwh56M/2F0jUnkSb8Mj0uz/spGDHIgkQCbLeV9xy7o9M
Uqs0zUk2+4fuOJaqAaA7w5VjYZJeblzb4+FS4D/IhWAb3gf90RYNnC9HkPl4ZDCvUpOAwNTaqNig
rFg8zHw5632mzv4nQMitsRu1Hu+CD5UH/SHx7QjmGJyBp51hlSMC+XpMZMDPIY+/yw5Q25gJG4Cc
6pjt30n5dd/7r+6VnJB47SAxR8ilVhrxuJ0MBOc+6EqYl68V8iefMbQ3QFGV3ygYbmNnMH33C17e
xORj3vBj5X0H2MZZ5nCJ8757ch4fb9bJdEULZkoJ52THUtUYzPjSjaXzI/PjKVbMk5b372jr1M5v
NkHt3cmja6HMhL36rC7BwU61KbAJgc5uEKXyPdN7yozBk2Yohogxm7S7NRlP0c+zr58mRcMHBRF6
VsfN6Po0adnbRQd6v0LCiPemj5uT4p8/8Zfz9qJGQV2LpuwsbKhhg3ZK/3yhRFVOeAKk2VIvz8rD
rNFKEdrmPPgsIlNDe6D77eNxenZqpakBLiA7xSb8Y1cNqTUO2hI3tSNqDcHlRJ9XWcKf/qE2Ul21
2qQDdQj/ByUaT86QDYHC32qLJ+HjC4OC+TvAvu8ddwErdQ1wvaMgMXjusq6ZcMyPFvu/A1tL9RQj
+3U9UMh1XemGfh/KuYzIJe6ahKxMe/hpTiq0ENq/YxSCrhqwl36NkUNP7yXsiqjGxkUUApVwQf0D
eMQu8Titg9sNpAtFsS9c8RRUsLA0LVvyVWn09yH1gn92resz/ZmH1tHnvQSkj0+cUbSpbpaiQGZc
Bq1cm04qvmMI/m24IgLa8jU6Vt7VR2LWLBqeWGSFGH+/m1r59A8ziB6xNk+4CjG8/AFY4aMK62uT
qtkPwk7jNLzJICiHz+QVtEeVMVQEJOmyRNaKAnY2q0eLf61oy+esmnCxrwm/vLrtCVTVpJQyXa+t
NRs6Tm6Nn77s5KvyfX79lBgiJMSjy3eBqsJAEoXioVthnDurboWHEgLUj0CVjJKHOyKBc89CxXrm
UZ+sOy6iW0JV5znlLQSH1KaxAJ9qPBnaSZHZV3U7WIBa0oMZiqVy+MrRvhBIHrFrclLLKvIieRad
n5wBUhBV0Akonuu9dNDaZ/9wLNMjVzaLcr+JY1ltPj9z7xa2wWhIZG8L3WrulypterbmxBeRpeAr
zOr80PJwquQG6V/zpe9NUZFW8bCGfO+vhRC3OcFx5xtOI9eJJklBDkB11dDLNebzkwcaoC9jFR7e
71xMe08zza1WhkTTsM7eFR8neJ5LEMPxb+DEcf5y/I9lXAwFG5q2o4B7L9pvsj6Ydwr9p3LPYo6y
Bp0gWbyalX91HtbUDotiz6gGb9kDiiHmU6IfLpivZs81sNGE31ksMPVwgVhZIOeOTM7lJlUD3o1k
QwOzQ5ewr4p7AbK+46oGqizGkmqnGQ0UTTjJ3RxPkcq/7xRanQP66vVfSMGgXiFlJ0GnhW4jyvzh
NkVFs+rQoVLODHjIdSQv2LWjlyGIXm9GU2PIDw/OhBrAdfmpwiH2MgCjd5+X381BoQNphd9qwbgo
UauYtETVKD60CJrLcU5EHUWYzeX/go3mMquLDl8WTUB39W3XGshmg575wNLRguvy8AjWo4scMoqO
Lh//T7ztCFEbL2AKXbK7puWnXyCEsNvYH0XaEcvIe3iAuIrEfq7XwIvTxGAMGRcUrwn8QqozXRua
LlMgzUebrk96UNFLHAZro9kLj3TC5jbKpph0Cea29CkOxOmG22tC7HxikkELzrYRhmrio4d3z84l
NCaMBRi9Pwn/oKgHqAizPUhBO8nf+tXXEU60v0z/01KyLSkZp3JjVnee7QyziG9bwf2VAH/eSIY7
Nv3oWWoor8128DasjTvIu4hVg9BDTBVuLBs8nrIiD8pmjAt+eF8XOmJsvs2YqtU/IrKvu6rA8Q0m
JWDqs3HYNYVf1MwIiRy5tgBFQIouFIvo7MO32yPPi3rsFzSLuk/PSrazBJp4ePVo9xbqX2OHfMdM
kRfjwDUE8Pvy4ggVUzrQaecWUIgHk8OhlHQu+hPEaUFsvSNBeyueIZ+gJxWSVxu6xXD8wd/J37B1
06aaEy2+Y0XWhn4C8pL5KCBhNhnkAvfH3B0jbbsa43Ly4w4CJ8IjpawZcTErB8Ppd+OgcOlFZPNi
4qhmVegZu65zomISwpfSIri0krFIWMOWtvQWn66M1SZ1YZn0GlYi/WXTOMPFvk1OXRH9aOMl5PCc
keAo+eI/I/rCQRxFMQP54Ny1kOGgTdeoqoZPNZMDulw+TXG9mijwz3kWJWlMkK15NVuGhALso8wo
0dskJ+rONU41E4EARTkDXkFaDM/fAyb79UI7gCwUSOKMuxmAQD+OeK4YaFXGJhimANgehy+byq4B
MF9PSAdAyqdyWpjxDh62zxtcQu6xIdcwWGV+nIIKaR0sEgTS/VQK+WdoclFuc9BPNhJUOJmH6UBG
CFjrcwQTzUUKbFfU6Rz8z8c8qGR07eSo12QsMqYSmJR8dEyK+Lne3o6lkB1qaS1TTZpAzgy1oDVe
VYIMIApSG4JBy8lxrxXaas7Rul0qtI69YfpUOdWhAr6+ZHMJpJ44hhEuLHRDnxg5UVgZrQRGJuLL
NkvygjYZgah5SqfoekAnkppIg4+TL1IwPBoaegviDDf/EZ7XevEgeY8bR+/7lhdkXurVY49g5s8j
ivGzUQyJ3qPB/TzQ8vL6vgNa7sOVNVHfpRhh6g9oWLHfpWIYcw7ysfocBtf7aWXv3AmHVnkXSScH
B3d9BWj6aOgTvIi8McQ3xJ5Y3L01O9znDGe+NuyFJPdjluijrXP8ryybCXoaom/lOTkBSOJcVZXH
/j8UyFqKVDB5uGeI6XS8OBvsTR29u/XpQ11990/eeeQ49fhSqNdXEq4c8dtBXxnzPJJ65zebya2t
WSskUbpbjSkDuNgYhKtEQnv9hKnkUFolPN1c691GX9RBiAdPlZahrGZ85aMFx5u/jyzoP57yvo65
geZSBvq03HQkgxOOfmf6MfLcjTuaz3IBJYUdSASngRjeh+VrWM7rHWwlDJveTSMPhgen4r/yH+mM
AdsUXSxt1jNeJISt2fQRGl9R/Bp/lQfp8uThQAGx01lDeKQKvGr8YwDY5vQx4U5sALNFQgQPoCJ0
flimf6FKQyZa/BdP6Y+nkUYQyWvRhamOjAIteEApHuV4UBTgaa6eZ7CCPYjfxfGwKEVH6Zb6/1Wc
mMJuxhfvT3qQEaagcBERszbFBDJPcxQbF+3sbn74L9QCIXZz19E7HAS2JgM+i5iW9X7h8pBJvsRG
hgGGzvx23GE+ONdGUBcSvS4TGuWI6pSYwli3UXpO/jDDdrl+QIcFCNDSUP1tmtTw9P+RQkgC0eXl
O8aBhHDBuM/7Gf9FPJUhAGLMBGh1K9TjnVgAvjw1zrUwDVcWWYx6TeEksWUw4TzB6+6FckEEnoQ4
0hDHsUaacy54Plc9wM7BRd3Lg8jQW8pYAkXH+pJUaXIOEddeufwSCUm2ABceiVy45uKy2MrgJDAV
2seEDhU2ulpL+cdI+kTy7nvrL96lYzIK+SLNQrjMIXWjqN4s5GCZg+bnILiBPBNEqjq0YCQhTmo7
BfGtxN9t5J9csdtF9cMxOMJwo/Ffns2nKOS3bGoax662SZeibCI1i0JWD5uZxomHGhuTexpIRn9G
48Q6EfVeXV9Yv+lOAn4ihFN2zlGHCXWqhcKffPFx4cLKA6hslwfxAgKQ+SFOwALdVSDeNKGbmSA3
F8smaDm/ppSr71lnxVo7+c4un8pGdg4AHu4DDTrXc0854g/6fuFA2R3KPKxiVzKt7BheWfk7OuCQ
11cybHuquqhJ+7OVuIoaVG6jb1++TBDWelrV37qgAYHhzSxugiyeXAPA9UFR9rAlgACMsNPK5wkT
Qv5GtWY695GGALYohitk2DGVheYNES4YF4VbboFDrWKn36t/yEyr9zSUAoiI0UKQhfW14NyftvMb
PrO/L8OT+rZWtOG2oADBfsFFLJbqWAIz5gfYCbdj/bmSk270/6zsAt5nB0IgwPZG+9511k88148l
Ejbl8kiOvJ9zLMgvfXnzXXf+2jOfJ24MrUhrCP7okJGrz/JkOKcAI9C0fJoeaiZt8WgvGTrzzPwv
XBnzFbekuwHUQnASRysdJ71CrQ+EWiPCkkPATU2nYGYlQieQ4gn7hj4ei4d8f3yhJZEvB39cHl7w
BK/1L1JZSyTtVrtCyrVez/1XNFydMb1wlZ5j19uINrnjz9dmpycEONq/d5OSeavLGKe1h0xyC7vE
6rdGO7B151MEuQNyln6JcBLiJiijed733M64ACrgEUcNXHEO3ckeNRsP7Apq8zWHlKu7ZqS4S6v5
Rkugt//Nq2i/ePY+0gobirgXbzvF4KiNP4Zo6zw3/JuuOwm41WSJXa1fhcZ1sC9RPreTJ1lnfi/S
JTKHO+5P24mMEV1YkMTvpt/61w2SaAOEaQSE2g6vvFRkqFFXf4bpzWLN617qPNHRwL2xLyWkinAy
wJ3lJXuM9wtoWs+4ITYd27kMOe5W5T214DOFy8JKtHl8z7C04GEvu/+9ZvwIj350i7939+nzDOSz
fxCXyOis6N7irrAY6jqEuNMkxP7pzrAuqSdIEF5Dj1iy6rdU7nv79YY9c9D6bVpbWs88jhjs8OzE
ys/tBw4u/dXjfXlBRf2HhRYkJEpRudRISrvEwkmMjrqGcReQgag3EFAZkAhIuExWuUIUcOabnao4
g/S3dnAWp3gDTGNmxv/ruts/gQdBHzL6sR/+NvU8RqXrvcSSZ/+h8XoSHSw8KA/QeRP6d+972UQx
uK9rYUfvGULpFm9379TA9ssQphj+4xGnblYWo/W6YdpmycAwJ+qNgoZnPsKi+Uul7RqAU1UO5gCv
hsm3i2wnz9N8VacwRqk5LZUgUhCTKaO44aWC/GjSFn5METUQEKrCnIUxl5mPxjEfQ3JAnXCAHOt2
NfxTOM2oMCOdEui1VjtdLQk/MXQRoEj91VNMxtsGUO37CLvZBB3JKbRXGJ6uQ902O5Z2f5vitxRn
7loCWFLrhmbaBIUw3Q7GF2P/8tfzc//Sr8+SdxxuPUVCQ8DCghYm+4/sScaUOfcVzYlf0WpBserF
XscINIqq6+OQsljlVN/p1kH3jc+J55JSYvNqX7P8TOSK3RulDDlJGhE7t7i00wY7uuIsHSF96KVI
yNWE4FQ0Bmb6MP/6Z7xnOi2Rgh4LtNYs7IwnZ8gk8ipGH9zEjokkjqDC6U9wWnFMsIX2bC7nmWBP
LdeAd9e1wL/twUvsGNvnY/nAv+dpgFm+m53Zx+1vGlHXmaLEl5YhhEH0h/ovVs/6M5ZtA3KL1ehU
ys28oux6pC7+6IOEa5McazhY/m7+1AvgIUB7QnlfSwQGR6Pp4LWaYHDwftaLUbI+LqioY8WOZ4W0
0+Y8KCs2SCQiQ3vpxAaNemphGaXv/9kFCOxSiEsIifjNWKMcs97A4RgOqHMP/dQixEtgARewDlCf
3FAixFzlaQ41q9mhFdwQyuBypCvbD5svXDQpoW9o89df6jC0DJXkKFyo7bxiOhQAT3wHfADwDqZ+
0R44i1BAHa7GfmnPmpDYOvP32iGmEiRVQW9QJtR3NwHtTQkG3IqkTgUf15AwqvYRgyZLWtwvbaZr
KGbHx+UZXDudtWCp52YSHlEf6hWhxlgcK7RotA2Kscl3i3IHR3sbxSYuTlii3L3P5/nHM/D4gKxg
u9MyA5dEygB4RN1MlL10iDBxXf3sFOTmXLHo3Krg2CozJS0lt36UxLyLqhKoziFZizNC9u9Sn5sE
Pv5x+JzY6pKcJoSVcPF0sZVL7qaVXKmhrGDX0hffqnyBUQaUtePsarqtW34HR4mYXsCnEFwDA1sw
4hDTuqI/zPABCHbW0Z+MaR1YQg2hLUvsDRe4zdOHWEoQ5ogWeM+gGUYW+G3sAj4BkkbY+oKxy5f0
YNcvPeuEc2hHuqgb3zmLEnwPwl8KzSha6djByytQ4DsUQpzcjgUeZTi0JTb07D1SnwJqWjN0zxI8
jXrrtfCYsZn/st2uubsbiVAWerzvNTGpm9SKAlJYxqJqhmD5kMRqxsDWZybt63r/59oxvoEpejwC
SULpRFDE8XtVKDhGu19uxTLHfDdAFwAcWx4qSMKQOJoKDORY28xt1OBwKIqZBuQ9xrwbuPAmE+Yk
rZMhi4Dd5CkBTpitRjRozRAPiQs0OOUNI1XX5q3WdaeMFJtoFpuWkgsa/s/Y0LVSo61CEG8IGhk2
2mmKNifRahwERM8NcJANuedN7qP6ZNyke+mid4kuXDMhKfzwbQix+WmVbvrgSvSbgpLv/Qfmt9lL
g6kaLem6Gl/ZmUmexwOfG+Zact0XmjdWhdP8s7YZNwA2TUQM93T5V0lWD38Peh5PRlAAqsRr9Cbb
aRzTgYRpWBpxW3dkIXr03fZdi/TOppt5z7RjYt/CxWDZKrJ7npLfIIfsHyygwp4wMK2dpXA9bF5y
Yl/v0eQPjcSYdGYBwo1HchtTHvy40d+8Q4Sy9aVVjhkhRNMYjDQvylf42hPiCGrlEMAoBiagQW3T
V4PUgIY3NGC4hHkV1IjPMFewm9JRvau+m/r1KdUqQgiE+UiA3H4QM1gzxOPzgGyf8i0U+pf7DNYJ
7GsR4MR+3W2NLNgXYqWiusxB+UTFKka6UJKzA1LOvkl5/9yR6Jwbq3CGtcLt1RFxDJxF76xyL5/R
HVssbsx/jgp2dVzxPoF8OzB1UEr5zTO9UKM6nuSDOSj7gAm3bCvlOz9TrJZrBqvkFjX7Qq7jeFqE
haYfsyI2AE4+HrTnqEOTbsouy66IXzGSz2c9zuxGBNx+tsg5qs30G5k00/3KyiGuiNhmUka5xuY1
ZqTmbV1c4GpNPg0DLgUhZ0FQEbamHtS60yI/y/7FxTkj4lo7Hzti9Oh3bhVjIyUT8CPyw1iDM8HC
i9Rc9E0zK3jsoovRNoD7A8j1YqxQOl9p6UxqlcvjVnSgXZlnjnbaUPOTaM02NK/lE3abOdGGG0X4
x7QXbhBFu7sKi/GlpDrwOu/tyD49K1DiW7bv0jou4iQrqZgPSro83yJcGsGCPjtzBVK3hTeoFDn6
XH95T6XNpjxvDOXpKSkWth6Y7fgSBgUVw+CQKjJPhzNwa6Tl60YsNCR0CJY502J2PgUBmr/pxg0K
lkjQzYIAGgobkXSprTpGsm7Ad14fKH/oxY8GAvf+q/MwhsuNpyvbvNX8C8621HNJ28GsZxH1KLyg
w+6VBgBU5maeN9xYuab+GMiLjvJ0OvKZCzSqD95UxwrtG9kLkurr3DoO5GGp99DnHIE5tuH1on1+
x2B7Ud63o/pOAlPaqxvCOwiafylaMt1fRnzQZMWT2CBeHBocs8DhJJmpTCdmVoxo0EF5+CrC1Ols
UaiAGbKhzfacbjH97GXp+lSOOlyG5Vnm5OOImOmKh7pHJongUKdjCsPJnGDgO6qprkLP9JnNaRjj
JLLomxVeDhKroOsZfuGSiimKCzPM6nPHL8P6VUQGXF0QejKI3Pkc7FQ73AM6ZPL1PT3U8qoLDqfG
1Xq6xV0UjScW68ps88HkGnDe+mI2/3MRG4y8bnVZPqAupnZb15QCIZ6AcmmyPTu6CVb0fU4C+TzM
gkhGPmS0JJ8H6sYDSRXSgzqJD1CxGAEhaRy6brXlA+5bGjM/OdlqngWRRH1RZKJUBEz/YoPO8rE5
3IglJs8racQFoSkxJU8Dbo222yxoRZ13k1se+nYOhsNyD3qhY4q6FhKe7eywW04soyy0MkmguXQN
rwhRd8shB1G+TTgqh27muKMiTeQF2V1vf5sLGnI18hZgfSukbBQGXz9QnrDQfDTR5Kw+d+6TXHet
fLMLCsJZ38COWc/NteOv1XKyanimorFF9wFnEomFag5Ud1JxonohvGNAKaV/FAaUZ496wcZjXoBM
L5zmST3kaULZdN3gti98xJef8c1eRox5rGyLQLwaAW/vVHiKbP4ID2Wuf0CQpunu/VrO7VCY3nRw
kTgKzOPVWfM9ppHN1/0SeHtMtSY4aqup/qtgxk+6RUy7Qgc8Ujwb5mkyqUvBtT33G+4Wdgi12ajf
3KxULInGYTFrAjp1sENGQFfsJcxhdpUkQQy4CyDLUAJQiz9aGIsLWe/Rfzy0uuH1mZfzh3SYRudj
LpBHWGPVcmF69I5eAZtt6sCIslPlpOY6ykz/mp/PTeCxTspPTeb5m/yAAXqnaRHEDiX2p4rZFsDl
99vUt7+FoIZARb6yywOYJsVi6HGsIEXoZaSdqo7fHtBHoJU3XNP5wb02cCsqBelhfvXcDa57+odU
KXfv/TUsYJA0JJ6xCc1zuSgWwhPluu937bIONpZDXcyQi2Nvxgnc9rjwyjV2CHEz24ev+JXTqM2m
DYIU8rTz+ae/YD3vW35U6yh/EUo/iT9x7taEc0LlNmbZRNzQFUQRGrfJ54dWuJjo1MT8nduO0EyX
oU8GvEIU7LIShHupKy41IwLxLGwJT05CTEZMJ6EQypzrhMx+1rYtfIYYnqmtbGDg5ozfhU76dEln
TnOZRqtQL4uT8KdwnUVdU1Qh9/STH1FyeG3hccwHk0y52BWBlwBvCNafnsB05ZGo++F2uOsXsqo2
DxvinrWqCFniXG7icX9f3E87uUVo3m/xNge0Vv2nDabBBh5VT6d4iqpO2nO/Al7Z4MF7k2MxUzkN
Fi8Qhw8TOt/rlqaR6OkWOC2aWGuSNkLxU9IMTbS8sCVW3T17Qh46jzT5WinH/NMUsIyPmpxPDrpy
FUhULCKJ2R11UvFs52kkLuYYs+cjoaSaFOMCnAJEtuNw2jFfJwtZkQM5rECJMOA7TeYHsw6aHHAc
YajgyW+NxxXVob4Sahis+pmgMUBw3oy+bpm2c/3NajbmTLQT9XO+aR3lfklsw6JhC68X0UvcjAaR
rs2ANr3z06DyTiA7qtyAdYvjo6GgvLa8TTnH67+NhAsboQYJ+AaBSRBLXSqOcL8jv2XNqzScw13r
f6JsxZ88ekd6thF+Gg2zAstsIDh/CzndN7kqnm/UTPPeoiNVuwyg8viUVptDd1znc10YjJVjYDFp
7czERkROPw4QqNhLclFx8rxrKU0XYPtKRR2sB+YonIbgEhacSzQIwf4EScZEbsZwcwZk9EUb2mHw
i5p29G1A8FgT8Vq3hvFKEAOtK8KWDPd8XSzS9EiMP/9I066+U/eoV/rkfhm6gwtQsY+iTrdXF7+z
oDhwaJp6bXmvVC0Lrb8Y5SOChH8xWi03lUKFYpZD+SPI3kYItXNZTksGSd2DsIitJt+llJV81xbg
sHqTNIhAy3zXPhzDsOzFrdYb71WsFyzLseM8SnNULPdicc0l2fOgt9x3ow6fB+6/mhcKth/YftLS
UA586rfoAhktEMmR3g1HzdriaVY625+LcZgqtMg64scnwKpgi7mn8dlm1xI45eGZQBYEfK0j+3vu
8pEhLwolOAhNHBkGUoY9GoeFRxD60PyjPKobwdTwpyhsDokZS75NW37FVcH0qdP8IDujtxD3KZhY
AMYgeOWoKU5uXG39tHSevqzW5Ou/jWFI+/4XplPCIxSNkbZZDBMBcpCSKpP75G6DbB14+NM8yMX6
XMHCP1mhKFQVKMBXCbtO7tp4GHYqgtYfp6xK8c6UkPcWl7Qy/Nn4AxqI5bjKM19vSK2EXk11h1bR
Df8fGA65GjyS/wfGYP9Kuto9gg8BqYn8V+gzhOgUmzXGxG27bjuc+C1uQeE1Oc1FQaEXz5VpI3mg
3R76cs8yL0WmbAvet3XlrFCdjH9B91l3rh43zkkbi6fPCrlb7IYdIYyo1ny/zpmFhOEQFZmQkaJD
MzwwYt3OolG0ZPAV2+ftLaqDXl6PLUCZ+7oCXIwbZ44GsNXmVE5FVkAlTM2invICyvKchKZj74C3
3M0ljDf7Yl2PYlSKta8/jrYjo2ADoUMnWJlzkpPlsxEnUEVsdjBPC2pgnNX0fvctnkL6x6aqwxso
ErHhZ6ZggJ54o3lO1HFiamKcHKSLXe3Hcn0xu2pb5X/PtoC/JOSckPTNiUYiTXD3G9evDeC4DcVA
EeAiYZ2lVjQFC0PyQ45mPQ6xSIlnxkW4+zMPT8g7RJX9Dskc4YTKvSSkkbUN/WFYQruSAUrjrtZN
kBb9e9lHfcgTvEvIdu7MYUYeC9T0u/YkC2e+o8JPd5V+tHW4yYbOH8YNbXxnJWwkyEAq4PbJdLsV
/acbb7Yly+XnC9h64wE0HsIZpLvRwvf0eiInilOwvadntnkvREQeL2Q6i4E/isuW6Z68kjgZW2rt
yOM7hPtDR2WJvhaoKLfq7oI1m24osXAfJ1hgJbpda9nXJLBCeR0u7cCwSHMQujV9jzicRp+EQhCv
yNNdlwzeieH9lht+UdX6digh3juJnlzPEoJIQ/BZt+MoC8/WYIaRgzvJzcyYnY1kAORE5/PRRMmT
1OLDGTpe5ybJyfmb8B6rS1TKEALaaRIA0GtEWvZZ9dlUX9NBPUp59yq3MQkA5TJLyjq4ZdnpyX+5
a7cgzhwqnT6TS1LXXziY0LZ5etzD10KOYI7HDisLvCvXEaqC0OoUc+migPdp7iMk+wW736O4hwqG
qZgRVwUy7QIVh3MdbT9yYUfysPRhDd0F3MlNu7KYpOaq6uZO4Tkjwqs/Tgpglz1tpsPt28lhxsm4
eNhqp6BWDl/dR+mr6xOsnAtDKOVS7Ef+P4MRYXAyucKW/lD7hB4OFeu/0ROAAbCVN4JcMNexQ49X
ocdgrJJt5KwBvV815yNSeITKfIS0jp+5IoNQuyo/39SGNtfD8ik0NnFWWIee2ZMwpgTtOPfFpKF0
d3Cu0aaCH0YvUSmGvOuk+uySdggJhRv7/ZuQ44UsHm6l/N72qNXTQAgs9T5Zld0k2Or11awR3KLT
4/RrMfz/fZ9mU1FH3FnNb4OzzFWx/wyKnlEOwOycOb9ygXfVAB9g/n2Xby42C/3/PUyN4I58rQA0
vo0YwYQwGk2KhJ4F8EDAuNz4weNwt6ubHpeTVnEZ91R00yTOB+VYSbWQpZEYRJKE/IEaR9/zNrFZ
oEwiFDhCAD0ykDcZNqqPkEhOKLqBo5u9OdJQ8nRzNOHM6lw6aPnURYeL68/2PUgSvL/YT2BMuqXJ
yKG1tojPy6e5RTtuAYgxWZL6I3PQYOct6Yky+gA72UL+RKSFcRxBE/iJshesQ4giCMUikX7RUrLm
58Nu5gaNWN2OETGaTM97hV/nmu7UgHWarSEL/pytWyv+d9Fpktqa5aRacm0IZF6d+V2rKdHvTxfX
4EqLVEoLwYZhGhErFjRjMj/sZjEcvue+E+Vik1NVnmJmkGvz5vnoBLMh/IVkuWt5+n5R4+rc4Wci
mFnNYSmglYYQbcXNkDIs52N0d+KvHjg62n2eNJ+MxJrwSZUcWvl+QHPBVA3tqb2EILHz13D+8Y73
bcCLvRdne55kBhh+HNq8kfh+FopC6YGxWZGfV3czPChynYlyz+TUWwXGZPR2lMtxuG4mXva2+H9A
PVu/fxVYqRI2IwA+jXVX35xbNNZxJOiSnQCI8o+tHpK3YYo7cb467KlRTAheR+/jF6tesqKdhfVS
QXNcb9pf1d9Oe1dmyDcflnG2JgT+8PEmWvRoKl4cQqiQQTaQsm3r1fzgSEaEKpE8A4BTurmCVFIh
vdynGUZ0x47YKcBZ5S8Tx48NiOtspoOBQWa8ZYX68oiv8iCNJkQWOHikT095FmAwCla5hqsr+O8z
mPuQPEVIyZKkNqUbG871Gy3MZXBAGAWkpoPNMYe8w90RHbJyUpBh9rAG+9bGc04Kz3DHUJud7g20
nRrd3uM9FPzuCD2U1OzhRj8oQdvdLZQlsUOZFxY7z94bUHGP5d0GVe+O9xTd0wYUl9vMLbMpGa7R
S1dhrKH5MlIZqam5UTn5gByiXhoMg4MknMBLotF4rmbZ2Vmj7KHZxTq8seRjy4Bm3BfVjkM3wgCi
/S3erjeMJsAnZDBKb18j02/2Wvn03VcvKc7dq3/+j1SKdLwYuDRxH7AHFCmlRGms0eUAlKTNxFiV
dTqbAaEOedfnh1wyOQ73SCL9hbD/4YobM/v32WZ1V/4i6HMAflTnEDm9SZt1fyI9e1EgWB7jtQ4e
u4T90HIDUDaQYOiJkyPeF7fvlcmiUvxgOZMj+c1+meeXCm7NvTbI4ei2PHxnTtzmnCN0wFw9XTmc
1ulXMje5jL+FQiQTtlQzRDxxUu0uPRYs8vdpPMoQZeMymvMJH6D2gmnVbuqKNSuXEqVWwzuds4AY
KQ6f3m53C+U0El6mSHSckcGC5hBimv8g1HcG1UQmROMpKDzxVjVZWXyuNVcsF5rksbuOjakfZ6K9
hU/fGzFM+3phZQn5ILoFFaADEK07jt3pDquu8eOtRU+4o0m9ErRaIk9QuL+wOMQ9j2Cbu5RhEZxe
+w9yPkIL8YHfMotf6FPLXYol/WDbu7Uuglp7HC5PY2U/EHxPIePZSkqIWYNllzVwhNPhn9JNbS9s
sExHzfuB7gi+Rfy33TeNaJjsrfAe6vkYCZx1Gq555Z48SqfIqYTwjnn0hsfocBaYn0IIJntC35ip
oLbIxlF6pED57d9iQ0v5UJk5eBQC7IWZh4W3+4SXkrt21tfiBsSM8Jy1do4kYBDT6EgdTf+O5WBA
CfTyGp5NLS1WMeny9x+PvScUXKbqUryYUFG96rkVsTxRhxhxrbkw27TdILe5+fuVZkiy5j1JyWpZ
G/0PHkawU36QtEIIdgjdlHXRfyeG3C3eyrwWNnlhWCEWlwHsem/OzpmNccMjDIsxGbNPjuAJ1vdc
KVBgCcOJ9NWGU70AOvHxM2YiCMQEQdY3jKg54lwNaqlKz16EQUHRfnVmg3cCwV3MCDLqilw7KVc1
S9R1J6t99K+dNt7kp/nzAFEdL4RvCf+VgpQ5J1Nm5tiICbkJOGb5Oxzz5OTepOW4ZxmJiR/Y11tE
Vl+nMlBODnX/G5B+krFgzDB3i50IfsbbSsBY8oF3Tvj2TALQ6hxrWU5UM6OP9JWR3Gg1sHt8Zpbg
KdvcJ78SMBA/V7WDvWmy/IIiH1NNOBtUyKzXpIUO0GSNR7BYOBNwOUaHa9lrUl06BAe6RgEv6Wdc
AzopiJIl/2YpjYJahh1iX2E3oM/Vw44BgA4yz1fiP2+K7VKbcYz8EbRn8BsP+S8sF9zxEd2tjbrI
zy/Fm+XMSoGdrtGFoEQYhigZhnaQ0NYUcj+wg8DZf64gcf3TkFYOP45nVnFiNNEWOChCbJLLEn2R
0aUR8zSiWtORwcqf02v81k+SaNy5IyoN6JGyoHbthJIn6ViZuKwbgpVmP9B22QJ21eksVIgtyE7q
gNGwouS1SpAprgYiTZ5mj4Ydr9557Lw9rrGSoRA/0Fy5/4zDYzkl/w/y7EqrMEGAIT9qkuu1/MHt
yxtZg6OkVMxQkPlXvq5jVQRL0+nk9YZkZ2vXve6wL6TAusZ2Cfdk2DSoPj3g8aAbJ1ttxqLIupSO
DLwo2VpdOUoXr5AlhE7LOiOWnE31GlyQ5mNFrGKdSImO+PhT2dLdvBFrZqIPQ/RvTPo4ncznPvvf
G/fEECj6jLKSYXkbBGMoe2oa8SDAs5FBKDps/1J9iiD+0vSUS8ahgT4Z+H/jYf/mH2XbxtzS4MaU
adBJV0mbyq1qpmlWdS/EGcnTgnGEjxzmgyz6rtDgebPySk4tzRtuH8+ADhcyTm0FOcEohURf2ZY8
GMXe4OoS9/ZoB8m3cz5j0yrnoJw5hOvg5y3fICZaD5yuBqqA24is/oe1cb/bHlzQssqB+UdasX8+
W2GY9DckN/B3vQflFgmeus7kxt2/KoiUy4eGSXQfX1tRSvVQAyJU74QDKOTpCgElrDtNbojWzRfx
ljWBEti+NhZBWjKU1Qttwvnv3s/llFQWDZtKnpTSH/64Vuo3RnxBSSQTqYgnd2qZ3qNTlPb73kzf
1jq6SJAtGjDqC/DKEE6pI13Qu+sQyyPjreQF/oefiCrhPT4bl2asTbsmremNtJmm+SzPRBlJP8fG
XdT1DjnhMUd1V5MpuQVpopNQDr+bHwlnopn+oQUTynKh/Ww0Bg7JDdjkl1T+VbFyM5O8Jsu2SvTF
ayDsciKKZtlWjjhSSdAkWUmzf/1lImsbkjYxYlRnL4xvw/uOnZiVng7Xvzgy077KvMf663x0dRHk
+GTgp7rdtMWznBRok5+5USyDnw/Qp1ufY+44+ON9O17h1clHb7n4crozMv/fJvRE0pYVq601rqc1
7nWQKe0qiWB7e9J1goNcdr6xzY0HuRKP9txTw+9QprEoLp/m9HDAccDqkPIrxqiuT9fXXFPY0Dht
rLUsILs4Gjv0hJ7sEQywzNNoCoJaH90XZoODJuAWRN0sk3OtaVXBTXwNEhGDkLqDbJVgLlVelG5h
GSM9oln+99ktSJoeL38J8FfjPFD5QPoIcFtKkkG0AN3CEwk1m1qaFWsSEbhnDuX5NmOI9YMkO9jZ
l4DZ5XmUym0gKAQnyfDNAl9gsNueUw+YR9iSdk2qMkjsxMYe/pY4rc50h/NbgIg02+ahUckS/vhh
7EzIk7bRG7hYuh8DEze2cNeWR7ziyHQ4HAhUq/pLbNJ4SPOEvtHDcEzcHdS8Ruar0NwjTVpRcrEI
5oZbTZ0c9UH3/KkJZ0Tno27UIV2eF6XYSj3ugCHMYcFX4Z/o6uUMIYOMkk7QviWDjqqTI32EcsAa
JcV3zZ+2LDUv5QHmh50E0d4nHZra6Lqz2M70rDDgkTjZCGXw4GBkGwOQEKMm+/UO3TZO7HSNUSnP
KHNsjmJPSexUdyZJEUrhfEoCcxsFKfKHd/Od4KEX+92OJP+UyAzKuKr96Gjnyt1YFoERZSbcRrwr
pKtOeTdSsIwCCHYkKUMtu5f+JHNznbjtyu5JQVKkUIcGw2QatAJK7qSsxhjrw63Y6mMVib8S534W
iBndEbgF1pk5nxsVjOw+SPSiPISHqzWdMF9BiQAcj8J2duHn9Cg7PYwGh7PehONFyIBWU6yHbIiu
QefETjdBX1hU7jCOA9UXVrkaMYjcPUe/v+4R0HOn9Xu3o3IHjeISjuVRawdS8bPV+tIxJqktN3vT
4rrri9GHWowarQ9g92pfSSgohUOCwT9WxI7eAdeQW9Mv1Px8CzcsSdKb/kDF/AafzOZ7acwaDwPc
hNQAEjZlP/hVBTIfs17G/z643KSDF/Bj9epZ1DqJaS/yUBXJkmhGBsQyISVnU4Q2KniN0chcwNuE
6gC8IgyxpeJhM+w6VIQwNAqMcq/Cdpnq1fr+9fIjU/jfboh0DClsUJ2o+kNGMnSiW6Tdd4rHFOTm
fJOBRY/Ba6zyykHA07JUo9VlLHnUl8ofP/pajfTyWmlreD19+ByRBfZr6xUMlwYwxwNABL3tOgWq
ahUuXCpEd9RMrh4QGYtTve4+MIyZqRhdvjc9JiDQEwTw1M9K9ee+2qugR8lYGKDXpYAOTTrCgiWg
Oj2B65lWinoT8TMZ6xC87s8XZKRxTSt5c0l7sZHbkKFWf4Iw4y+iPRIumcMp/TvoQ5E0PFM7vAqi
WQRmFjOnKSWoOzbS6jDtLwOo1/ox+uxaqDYWT9X83eqOpg/ZJ/REkL3HPacrggTPDiIQKCCA1/uJ
TVZnxTSSUUlaR5UT812/FZ1cOKIXKGETJ6/3JvLxw0M+yw/SK6Ty3wrm6sJKT6IL7kZMMxGfw4m3
KDFPyLStP3CFOkv4SXRReJ4RVhatyXGA63KTxIFQ2oyBMYH81gENXJEc7THIsBihHuxFBAqj1zZt
bhm6ePXQ/ZtQKHW3ZsmKuQlDkHmY6Aqf33piSRlGoUylNgcIkQ0WdK2MJvjw323UVC/KhgA9Grk9
95YGO7TiSr7fAMcMXFLjX9cnOh+2mSpCsUOPgMmBSjPUW6TTHwJY944WiVix7Rfx1INyat6NBb0T
rKCRDc0Z0a0U+vIOyvDth5BxeOVrrOCjfpijq5RCrBJRUYiVdNgni7OLiSOvu3HvHtxO0c9gtxM+
8cEMat7MQqFkPG2SXl+ceMi4MEUQxUlKrUbpwYrx3+Ss5aOo/txx1jWRq3CQ71TpPhDRxuKR+w5V
AG9AHSwJCS7Jhr+YawcTnwkvnN2Mcx444t2wwhELw46y52oKAcf5E+Yo2jWfxVfpNL2I/VQbXb1k
jv24p3zxcROp8ycrxBEtJPO4uMx+1sdoJZ796puIXcu+1hXnKI/hL2MoC2pHbTRbDYVV204UYcSt
+LAyORl0CHlsRTq/rJfoFjCVlCrbteu/ps1k4rSBM2BKSA3SILAZwHQ0AkE9nm0yyFRXrJNHr3bN
IkH6xeln3yDpglDqFhOI49J3ZODvMItVo7ZaTqZ7bK+KFryPgACTgy/wZV+RUXEEaY/CTzxHIUgO
sFc9qjSp5Ix6Rb5JC28RsjiWZzseCsLRewYmRHm7eqNkEQqaT4S4idWfONT2uSDYYi9JADJ/iGQR
www8rfi7sn53nLZKYTYvCd8oPRmYRflNBOfOsso9g3Gh6h68pGVvw++af9KPlYm2MroDQ920X5Kv
isbG+Q9lpgqO6z+R/cF6MADxc7eT5FYVMA7JV7qwtN+8/cQ9cRc0m1v0CnHsEdGGHWCUEfTNL9sx
eTKRUwiH4Kd0VKsZKH3tf7cYVB22ZQgfQqRVc5iKCML67q4Cq53r2T7W74rKTG/vSvAjQ7wOaOsp
/o7NHSN5UBw/4M0ciyYWU0tP2gsnFzuZZqElCP63dL4waItjjaWejkQftG0Toax6h/Ld0o1hUYoV
uM/vf2484GxngBWONB2Sq+A/rzY5lqUSBSc4pwZ2o7sJ3Avnd41qeVja4RhJUdX2+43AJYwuJijE
CUIp3Wpm9LpA/EZSapp/oCZ5WQGRXDb63XQEi5vzfR+8KLg0JBHjg2WjUCCNEtweHzig2oPsqMY8
if9b+As0WRCHVzI3JlSpxAaml4O82NhlVpfJone+T5NPufy2JqZHsArsPZAvCBlz9YVQbey5YvXk
DhbLHvyFqefO9jCb0SDIgc7hBfjGAJ/tpxj2jRCGE2Wehqeh3vhQH5MEz8Gk6c8PApkKquF4hcT4
Bbhoq6WghgaZ43N7jT7cSFmgaS/OSkBsweXC5+YTjIr6lcBiEjiU3+TIYuF+oT/aQHy96BwfX1r5
QMLkOujBG0iZdeXa8g1Y6Fyez/eXJuRxajWkcGn3ObOgOAJ+TxVVl64SMaPiZvZoaxBCn/ifO9Ez
Cj7jgIk3EccQxsy6sQ1q3bP5nwMvqpOQYApR0DmticMr3eKig068ApXyAsYd9BD2Fpa/NxXuANaP
zbq5J2SgorK8UhfPGcdSYjI5bRimqjb7VuJrmXBEyzecbct4f5LvktDsMke39KbuEi4EdftCMI84
6VktxgSn356ShjTXLJ3e5QrXu7dZoye8e7CkXdt6R2rsPqmLAq3yJh4A4+5P7yp3GJjcRdEA8c3i
ysjrovpHzpyIjAUbTRA6P2Jxr/APr05jPJ+s2fXf1NLcbLQzDjUn++lJCntri3/k9MfGcRirXgX/
k6NYesrp/FdFub0L6hNgANBonwrkIq4LXsTRggHQ68Zdnws3SUGZu8WZbpH8Gw19iQaWtL/rxbDc
a995irRbet29l4Y4siNxwI51zqwYTr3I5TNAQ/2Un4NYC7ceRgP7nM+EI4E1BDluP6KMMw6rhYWk
rougDnPMt+sKcPcDwDGnoDd95wjAJN0w1eeAKbWkUyFmxWx/9Gn2YOb07jzIQSEgLYhGC47zVX1D
taSdbl0BV2tYilnlnt+roLcwWEHuzpB5JHrFNYc+SJsrWvqGhpmf9V23AL0Sk43VUwnvgTWQk3ap
En4+15naSfbvEZ6c5UbwINi8ykpsMwUizNy0mQzAa1ogyuUqhlohft61k6DU3D0aJ8odUFx9AWYm
05uzOq3TpfC+LEiYs1nJtyqE2y1RfbqgmA0QG/2cRtvpDYGoHmkrc3/EVX/bhDCKZ6hvPpr116xH
KYxafjqz4Gi52L2eQnmdT0oe+BL6TllyVkIxLCyt/lAU9Xz2VvWNX5Mx+68Ar/V1UCP6+5L+OGbh
2h+hNhhCEZRiTklmh17uyfxrEMomd/wX0oNPGn+54E1I2JV2WGDfd1U/2DL5EI4lE8sdnVYYoJCs
FAOrPODRVAonCSfDHpD/M0B9YhLntKj928P3BHosRWuGArsPowYgfuV+qjU1AtMbYn26tPS3R5NC
08zMM8JrHdfqONMAcAHNc8Pc52nEIKxSzhFSqlw+9zxcs4mqHrH8RHVgoDbTFoafm1jbWCWZAu2V
a7kax0PqbcIUWG5fXQdXU4n9fN8RvzCE0ryPCIQZEZK/pXrPDKfGsRIh3dyEQBhqBBdBvFiwOkUr
jQqIFiC1t9g4xPam6qfgCwr2FescP3BS2KCjbog6Jb12VBX9D7GkWfJ2wHc4Mp1Vwqw0SkZ/9PXi
LN9pLPAUMLxKHQ6+MA8bhfoVBJiMc+PpJ7tYnbZ37TYA0Y+q/JVj34mRCy4BHR7jJZPdcMxhQNJK
sDLui8gbQd4aNHbN5JTaoVNedNoBcSqRWSlNoxWoNwDkJPY1TwnUkrUZfIQHjziceySL+qo59318
djzLorbGZbHHpm61g010TJUIpUEKXabNg+Wh8VtCHJDTx0FoWp3zATRIDx7r+VFoEkOrYCn6HZ6o
jfv+Ks6I8NZLw9oTeZsCaDc35sUjyxi3TVJm9ng0750gQv8hJn3o0RFi0ohqsDMXuIqMb0vlrJHO
rhJHyZ5TWkgzQULQXI1gxQQEveiiu8mB6Q9O4pKxQEdXjlV2e/c9bikm9/NooNcl6+vL6WjPbB86
GBdSSF27ve3ytWF5izy2y7endmW3Cshe4y6/DKB1BMBXkAfzfDhXGbnPgljfPA9h2+VyHYEHeK74
r1HMJA0R9kqWYcmDBh7SJnmA0iTKZNdtt5x9EbtJpWyQbog8eBA9M0PvVFyzx6YXhxu8Mdp9LZe8
BjkGp3ee4W8CnyD04oLGwamE9grpvB49Vs3WxL+c809gMXtW5b9AVGUX9c95UQRsc8OUyd+OpNVu
Qk1fc2kD8kEXVykO//HdpUo0F3sucTZQgF76LwmAtErX9Oqrst+1IRT13y5EbrNSJ1eXWdW58AKi
VqQh3rkuanpoi3Tr2ZTv7mubajx5ETl36IFAVhyPfSzK+hZ9mSs9Yr/1tSX3mTLmLeFof/gn94VE
0HjGvC9Uf0y5VZC7wYzgr0KlWEOyL4mriNFn2HisXa9yNPpSHdJ/Mojz36g32m0p3g3M8awEtfHm
j+6RC4KV/6Vpk5w1e8KMoj+0JvisqZf+Cg3ZemoxT8pGdjkBdoYFo45yEJAmFpGuFl29bMRX7jHw
jkhXB43FetlTZPhLb9GbUxp3fl6R+8LU3bjQsuS/DECheyNIq98r4eYFeM1iFmaDIfHf5QdvDKXn
D4DiVISnUeMwyaB0Jxy+efTaniX/qcfSgRkv30WUSOaA8P7gHhceMYNP4S3i4Lsjj1M0yPjJo0iP
rLl3gFdWGdboo7i1eMV22VnOlMoHoMiUzpoFpWlEikEyDs/4mxMNmJx/3SPdnx9HYsBnrxgvIth1
URuo/BX2wV9W+xVHXcRiMinKuu8iGlDtQtgNt7oTWDgIDPNq/jvrQWSvoopnWrY6xwHdufzBeFTN
BixqXa4DoaOXQwlcBWiA+Ke4FRBn9hhQmZl0E0Jr17MQuwxWnpfF5CHAz6YbTt2aQ1KwxZrApnWa
ycjkYvbdOaNmAA7kJJzYgg70KJT0K4C3N1cSv+RbOvvQifljmAGsqZ8fO3acbORsTzR3cEP8kIQ4
tyHsP+loGfS9ajqfys4D5fsCYX3PNqBWdD8o0ejBGW1cOPG2ysPNn/hgX+m2szzuUn+7v4kLwrHl
3d9FLZ2QoaBeyMgEsttcverbxnsEB7Jl1hWtsFgold68tN1S2Y9qyC9eREnuHXDu3FDX20EPsXFL
FCruAklHOoZA0Ag06e4n6kCqCq85AYdnXge11ul+wMvUeH8iZWgOy6EOkvFt0+YkF2GEMmeanfjl
n0UsZcvLT49hTBzIsCJT1vW7H/j6K61w/g92Q5GO1v6a+43a7h8KmlsxNIn7GRC3SfgPhN8v9LY6
No2/p73SSG2NTrk9TxeI9ZiX4Mdajb3nSYekSb1j9pRTW55KprYCAoVv/EXLmCs87wPfZXw3f5uI
H8irDsU2qiEtu3RJO07rZLjCPo5Iyzz4qG4Hf2IKh1f01H3a2IpbsE+ALJ4uB/PdJLcV0wUGOEEp
XxB7Zo5vXpUmcnFZ6Zr94vhefFVfwkpetmzioUtNbiojaImvjppOWQSSyRqfOQiUGdt99ApmeSzX
AJ+0mFcJt1Fxb6re3tG5NKXpWTLYDISEG/qhXNB/DlQ0GbkNqPKXQOYQBoNiS7nTKKF3ZQwpU5mi
AQi2MY4zjMyj/DQORbTCn0YPu+oR3QfivEFwJHu3K8h+BP85ZpDc7fZCPxHekNKLJVCk/dqUZLTv
rCJ9x819c/Vc9PgsxRO1LGObL304oI5GPSX7HRgwoVpo6qxbSfKBthaJiK6OWhyFk7+jKF2EIjdF
mCmUWe++AQMcFUX1zmhXFo4lXZoe0RqXC7FWgr27jA+o8BAgrK6JpTAm4vUW4ZyebCgJ9iiPONPg
WAvE8we51Ihk64KgXtUm1XNVwj8958TdXiaxiooMElIy+1U08k6Gcp+dqCMC46VkdpTsh1hLtbNV
A3O0xHtDycAj2wj6tTkHzeJZjyjQ9jCJq7MAUvN6kgdXj5ciQrmpG8meqP/ZAGYDCMFoyLBmbJtd
tor4l1l87q6LCN/BIjr9G1Qo0+qKnHv7eM/aUVkncvAmWWIDMdfND88PkeCiPx+TraELLUjk4iAM
43v7J8NhHJBeZ08eqxOOswSE4YfCx0zlIY3IGimWiCrCFhZ8oF1I74UomBvIA9WBOFkL7Ld+v+Hr
EbkYDww1W5NU5hI74zJtzEyOc9C8jeZqRVLvgV/j4E4TWTKldeU2XIuG3fxakuT4qXl2dJf2KX4y
NfAsNutwqk7bb7tr1lA3BoJhqDQjxjWTzBwTXkc1j6WRBF1NRTlrFz2sVk90GubNvPSvB1WEaVLs
8mRisF2KzkI1yjwCvxetuE5rE6RItlWO1fgAw+0STK7XwADXi5MTzYofG8hbVIoUagxo6gCX02Vj
KPSnVk8l/DPyPiDdSbqVqtC3kcUOvl4c0tFoqktTzaoJoee2ORnyA7xT8gIg1zvAkzONZAEDosRg
RhCLg+/HiMkFi/VGpp9xzu9RPFGwzN2JIandw3MxWz5yWcFjBqOOPytQrD+8+L784v4QKM147q9U
17NzUZBafulVkuUY+9SHC9VEJ+qqW/z3CGCoN/Ns8G/c4Qjsu+DOHpqKjoghpl/8MDxSFVeFFJCk
YmUjQgxenlIwsmLHXVzhXWSsvFtqNsUSncc9BVDpy0f6MHGJ/YYZbylo2BBVSZJy+7fH9zupyhEN
vtkNcFbA/s5GWY4Wol2Eefgp80ftOQiCX0SV1X4QkBdwaiXYbpGKzrp4UQYZsIX8Q+dq+9ZzApDT
jPs/6or048vF2E8/ezfiP0d24X/8jHAFslSJPJFj82NoPVpN4RhzqNeL8/CFD4z3t6MORJsjmA43
fOldsnZTyhoYtr96JhroHtWimQpb6I7kvNfD6x4xlg5uUdq+kfvB4qAx2TETHhb5fvglDqEVGybR
o1cTEchfA7NobAMMz5/yv1OaAeTT40HQ64p/REy9Wc3AUoWoAmAuUrbT3DZtDGXFD48u6xWBuEyk
LICLKcrJT7xLyDtXGBCVInjPYOIyLwejdRTrY0kvzZmc+lZBWyv9oY8oHOnrwfN5Gimwiu5UHSx8
vZLdLDMX2NztK+2YlIZqYJBPof1tvlOHnx84MINBs9VJHYzz7+gt2aXxjEYH5sSCy3w2gA8W6Km+
U0MxITHI4g9DV9+Rn8Vvf5vndcbBt1XsifE0TdSp8/HJs+ndo6jx2HQRdzIwnTB3Io0QZv0NsU8d
6pffIfPwcIrYujaYXpoC9KF0E9ZGQnn1Y+Ky5Doix9VX37kF6Y5vHEbwVbf7fqxQwkMoE5xuvX2r
uRSuStwOnUeIql9v1Ddsgp1NNhZSfzuCoX194niokehmyu5O79qLI7xmglApT0uqdnYxWXArfFHt
RT89REUIAEGtYqN2ZXhceKrwFyiTTywa/EUTKE5Z5AxeDQyPfqg3I9Ou5n0OINXOTqTM3Y1FrL2s
9RqfQ6JK4MgHNAQ8zZ8TglVkpe05Zn2MYpsTcDL6+SgH5fxRcNdoV+VYpYdgDzI2K/R8eqzzv5ER
bw1lNyz1hP0g4IiZn/eczBxdETUCb8ouR3yMwCTGRpSgpuZkjuVYiVze6Fgmvf6aIVV8ah6eAqSx
9EwRiTryCsDNnGBzk3m/me3D9TtjTNtAm6KO0bfUg+xl0NN0O3RtrEna7o67jsmY0qgWyhRj7t2j
zDtUyqL7rXxj0lI2le9rF07UNZCgJ9dlTYLoFH8MR2Kv7YPvZoyx/YAJ8TBhOckCQi7lLo3grThD
Pwm0yShs+fFUJjyAxCwR3fjJWzRS255yhQBEryXeK9TTQnAk5oW1Ib0psc/ysv30/NhlZdZAGCEW
c5B5CidayIqueDWfR8ayF9KJgZbWTTQ+w3KIm0FaxjVaf+kLa1RnRHOsxq34CEmosRQ9E8HgYn8b
doptW8fiLBp+YXQ8RKCVtGziZoA5mE6paDjT0sqtpQ5dOdPM5AX99AhGqQovyU8kkNzo3+x4KHE0
fvomwcNkBMc1efMrySYE2p+ducjPtnlHJtuuqXV2lseUE45vPVnr7G1v+xHaJhi8hh9IAMr6z7En
ffT30VpLkdk/BZQBNNeloEV0MDEkL8BBr09FL4XAT2oLO85GAurz0N60T+dQ7UUpDKJ16jQwW+iq
5YBcaUsCH9O6soG1ILaDMA2Owo4qBHXV9io87aBoxr0hxUucCV1JH5tn/NVhd41tKA5XBKcNVx4N
zcgq5/3jJeR1W+7dk3DIgl4BufdwPYpiHVnhKF9qEcu7l/TMgcVu3C8VzR1O8RsyUbIJKEaqCc1b
b2L9utFztciOtjzZzjJtCRTfKAcMMLj40lHgWPPS/WszzhisxDDVx6lLzH6Pw6IwfTvBXj4sABeR
2CXqKTJd+SLxjYCN/8cUXtcHTIlIBK4nu2XhxAMU4/C0PsH+xJ0waUp5H1x+56cd3CzjW1bn9hlB
Mer0YSaJDZgNGMS/cKNs4EuBsqfZECEpIFK+fHXBAB3zkD6avNXeV53DneOmka6p6wPip/OhN6gV
QHxsXPgtKqP0sww/QCXTgDb5SP+f1JNon70HuybLBeo/xaJ8VuKtBWs8tMfv6AVj92YWM1xlHFG5
wETdYlvkbQ+mN2pbkfOcXav2Q0cuJ2HkcWklmygfzBVnsSRARMeNlnAJkb/r934QAjMbtQDwB2dc
WYNTqYQogQlNz5BeZogLlJ88iCtHlJjsiwb3hSKDBSbuHZyLcI2Y90vzJ4acZuTtp1amW5EOCaNV
YXU75oRc/Sk/0+QIdyWt1AvDiTIsSTj9I5hgNBtBVVrhs3MtwfjnJn6iDQ+SgTwxhn7Y8ebzN6+g
t0F4f7gjBnK4fMqWBzdHFlU/DdsOnQdpM2G2f9ofZ028YCAE5uFLv6Ar0/ux6PgdegEl60VLn7ra
+qllgfki2RVY1e7wt5QAj3hQcW12s5umAKqP9LI8npnErdyVxTn0lpAATuDHoKrYDdRS1NoIt/DZ
uii3mFQE3RuFCLI52ccXYcaqB0tb2VvPm7ZgE2E8uXejSbj5CgnfVR6D5sslZnjpbCDl3Kwx4SqS
HRe3qeDDNV6D9K8CTe8NvkboagfDqdqRPqh7H8cBoUKDiut1gnHwm8b5/L3ybKAeu4ajdWFDXigz
z7YfHo3/Wk2GkHFhybB6fCIaxIk7If0Z2R0ZF9AREqyd8+dA+UggzQddxOKmfTyH62B5N7z3rQDj
2nunrNeEt8XieXbdu6QOVvs/Lq3YVm1he+PWJUtBDBB0NSfGPt6iJyKl9eWshOWr4QfHzloBalxG
9SrRdDgTI9OzrqT3XITe9fiLrHgpi24vs4vVT5Uws2ffjJR7L0JLDqK6rzhe+eg6NkEnSmoRIvV5
niVaDSAOW5WEUTSzY6SlTIPG6rhkJCYdxJPiOzBcgWyV5Wjp0GPRZbBOOw2KyliGF0ArRLySPa24
ZU7XurYbERIP1lz42AclwIxBqO2aOgY3rzs3nd77o2Uv54wmzlxhXSNEblgg2/u0cupWZIvsgEGy
qjK0/tQR+2IEBF6iYeKym04AVsn9Zg633lc38qOrHbQYYmWW5597NSW+xhhmWxgdJX2cU6fIEqTY
v4GzKYjcsjOiTTjZ1SHpFbGDVvzUXX+KBwU1Y9o5QZFixnetTtUZAe8LZQLYE4/t3lvwK05o7k6m
iycKNHOok3pCC5rGzzvDIMcZYv+LFWBSxuJmlhB75KTE29Ux5xCJN7FE7QYKNy6XPdWrDuc4fZk6
u0M3mtye3f5a/2X+IbJ8QxsiV5DpsQY9uiKcJ7GeLYsDw1gatYjaZiffHuqwcL/fMjEUCdG4djPz
TsxpTxwQFodmGQ/OQKgK/LPSu5mCfxCvRJokmEFDlycI1PNoqfDf1s1gjRv6ccpUeip+ekcMkG12
ZrQT3XfopQfaPxCQZp6TDzLBVFKhI2XhARdYe8AQF2Y8SexpkP/YQdKNw0ZIE+Qalc4TT8MhlJFe
a7DIbYT4DD0DNyXMp7QaMP/zjl/6xhPLakU9R7fIS/9Y/mB3jjjdiGpCwvO2AHj2/x/jMcaxLcrD
P6ix2abOoOnWTTwfcZpaUpqSyKIm/KIeH+k06TxmoKOb9bWFf+Bf++18bBbLgBWd8ehSclESmJRt
DO1w/vj05gbMNSrB8HfA2/MGVn+v1mrBBAqCm469nC5tkfGP4sI7eg8NOypRKtQ0TLilLKVVUGRj
UQlS1PBnCDZEG/w+R88x1qGgLZU/BcLf3aweA9aAh8F2osAb6ZlxSLwMRenPmgoPPlqimKhVfXEI
dUGUPjG4YEV4R+Fd4xo1EuJiBw31cQftRZ6u13Vze7+pOvFEceziU1Iw9zR8lHazrpi02tHYETyr
qCJZoE+jswXku/Nab/NnYOjbzwjflWayawjKC4AtB0bel/xmBSnfnSPhOql2ReCAUpdHKgVahB0V
tXs9PUkveUHlly5KmePEW0SDNZ86xj1k1/gUsL31ZCaXrSenkKDUcx2f+9DJ6ZUjscBa0Ah1oYg6
cRNiYxtnqmi67fg9b1K4+tsEFx8Gt3v7o8s/Z2rqQwN1U0027KTbpo/+PTGgfeSTbZsK1nytBe4X
SClzKBLFhcinGQO9oo/54rucJOVlE8daGpI0jUHwIjE+Gm3x4+NssX3JcdIFXKHb40qoRRwOROLW
bYV2p3jK2IegQmahHhkVlxbhNTtnFHkgQujN3de6wpJxzCTJn80mQN/UopxIgFtJW4lzgldtZHwk
QoxeqLxKysfawqducuT5V8a37yaK2qskIInZduvmIRpJFwYikVwTYw6evu0xoK/YpTCVfrV4D+Id
jx4FdJikCjVyWRjAeF9ulJCEveCfIpK8Dj8NFsT9caj5H2SfWS3oU8e91TOWFCMcDYbPlTDj0pl+
l+8xPHR7WKX7rrMxHbbsB/LHqc6C0uLoJFdSMwzO1m7NmDO6jxBeaREoN3kI97ew9QDxWWqAOF1b
GmVnT06/ZHgmA0QjOjoyJrzISTQv533lID9e68os9LKSUeTG6N/ps5D3O0ai0SI6ArCTASmKlVeC
amiTwDVzBhp590hiyFLR1YDHhCn10TK704RisJaXgI9DzbC8mSDGuM72idXmy8r/VsD9Dwdi18EW
PKQepWD8Os+SrYDUW8ClzLQIOisqGWw66b874YUys6kmVfID26N4nCvpverKCcMMJaYSpDhrvVjm
7CAnLx6REp1cHLt5ZJNuB80ZHUE5aljzngVBkOjNyb5I5S2Vn48guWYoCtkr/NIk85yKlr4u1AI/
9++EI73Kh9CSKUtrQD/yPOyExvVfukPVMgjyQTkgnjAR4yx7tFEskvtITGVIbyOUE9Lk6eDbtg75
LcgBEqUwY89Dwhp0z696M8sfR5CVIUYzYhyxn/zGsGKMqcPXljU620YqjOZU3KLZKHRBuw8hcGaZ
q73NQiRWMGxCFWLbnCRvW++wywLOM2WIafhMuzWOEgQkQ6gV9eUfzn3lwNE3S4DXkDmbEvoyffIl
KIjNV9pAApO5A0gNZN2/XFwdb29nN950lIpWyUpj862Yr16hk1wwYXa+s+aDC6M1hlR6ahc4+a25
1j4LRHRcduCN+1Zxlcbi1/6gACDwYienPQuEMlu2w3I7oGfWoOjtEs3M620s70Dk+TJ9se72OaM2
TMnifoQcIekhOnxLQAQdLFpKpMaV5dcnXDvDS+OjYkOO2HOkhM8PSOVkyIIv1NDpsvFzoxYwg5W7
t7Z6ycOg1aENYZg6YAGVQrLvsmOkioiO5JjlcZIqSTD0btt8Dtu9hTcAgAd5M1oyVYZf6XzCch79
iZZ6q7VRN6WK1fwxpe09Gj4tTXjEN6lV1uskbmOOd9YZwb7XaKioMH0tym2NWeGj1fU7mJC2HCjC
h/OnPyD6ZegAC8ekTw0rBcXI3tDzXbraVWXpze4QgYsiFLFDTr6ugitBeOcWO2g+fN8TS0OpddzE
9we2n4oyVvPd88POftFQS3WzCXdbr9AvFvbfHKWxRf/e1QB/k8X1AbzstU8FDwA1y0PRiu4HFgDy
gJGJmJqlv7scKLx/gegilHJg5xz9BiOgryN++i2YtOxzIsThbOp+oGb9obScbuICaBD13uUA7pqv
XAGEjji8ASrTw0P0mQQ5PgW1no4uYJ16O2i3Tv7Z2vwpq2zy54X1ODtrnUkyPXRmSZBw0x6LYH1V
ACurJl9xbGUBjoql/WUsvhhKuKUhVa3IqruUyS4klawSalCdikRsTvBvUCHeAnJehY+7hDlNrEV2
0Rhoaw/JgQegFdmYE7IXJCKV3oWtP1h6ddyNVWk24fMthjPI+tCOmdUCweVctzgYLznts1/1FByd
/tAadDzz6EShGu87D2RNledmm9ZUPcd0UKvA5mCt2Q9WSJFzeEqh83ftIbgLxi+IAOLEGuzNr6DZ
05p6RWZOGjEivfh9FhNZPeJaNDHffqSZXeUA38RCxGI2aXISJ0zAVxyj0L84fC+Dy0QX6W/yEfC2
R+6M73kdfMKNPb3f3vsWkTWYvM0tMmgrKp5IQVKHnh4/poOmGcX4mjBTmrVN8aboCHt9OJg+D8px
wPpzj9YkC4+oPT+LxpyGs+h9QCjE6xDHXgZ/Z4LOXA6UISd/X1SFWylAFEfrvGN3E1AyEtwQ3U2i
U923MoX9Mj+pGBt9s+XjZkpUtYKTTcJVynUTmevJRqe9bNTT5/A9WM/DyPXyT7PXQOKSjP5u+Cu4
Gybw1qCkAqN2u/xauxvbPQAjfXc3bO04Yes6tT16HpMUuz+Nc5egplPqMSccOtXSol0akt1andsn
g5sA3qyqnC8PQLHtzjXnzOsq/nIMZEIB9xrWMNY7kxoNW3Tk5x/9eqdvrP+PJZ4RSGdN8PQKx1kX
zX5TPT0WFo2zU+VcuHLIfpAHDo+PcFKJO6Ck8NZSfGFy2RVGzzKk/LnR/EMLNz+YliHNvSJ4/maQ
hJ4kqG5F9x8fDfcRvPNi2kbhcDOoZPXAdWO4QJTm4FWM0LOdgtgEshoTW4jAkBQpLKMCqlwAiT7c
ZwtFZvJ9xtVUQiyaSzpn/RFeRRKj4lpEMr0YN/GbJb4VI7Sb6QFJE/Yxbncjs3GHVfN5XndbKBoC
9UNUrqJjHam2LKDlqYNm0o6eGE7s/ckDReRTb9BHRlFjZfAdhFcmtdDkJT/qxE48oziZqlRcD7NB
txgJwIgnBE8/rozKMx8yPJ8ofuqVVGi9P922kqp8iTaFZZ6qXk5UItdjW9ojI+1VSwnExOPjEGtl
vfQLqY47g2kCvG8oMZ/7wM4AHWK5U2vw70KrOY4KSAAanfVJ+1t7ldHXxH2bkPj2rb5hieGvm/4v
ykWnP8uT7M2odLlwy3pvytQxNbaQm/lE+N/r6+YmbOIy00SmWC7CqATBngToZULRSxJ9wMABc30T
iVTLfDaQrJ8/WrIiI1Z8rkR+gbMiyi5e3lG2W0qDZgCIIlCbfmLeXsJV+GnnYCzunXD6sT7Vuhcb
SPSkbYJuVU1pmOBDKUY/aZ91pOUnP0f5DAimVSrY3A1XnimXLaEQ+aj6hg8Q4YKrjSoAxtgGrq2w
v3vobREDDVk9x7ytF4wbulV5TQJMAUx/X5qCvKneKfqak6SWN+kwyDIaPiUuQaWxArstRY3YwI1o
nPug/4qbf8FEEOMJNbT3vN2ukp+CtpfhSd5iV/SJEVm4VujLPeKFQNrnuCGlQ4plm47f0YdmLyzs
+hWCGk6RIlgUhqG2vd25+1HsHPJGBQLJwo/E4tpMcY705OMWtKynkXUxpWZucQ8hjUo8oCiI3Rg9
vPVcXdsy3OnUQ4Vs+TQixN5ocg7oXmmVG3fiJvw8UK1Lsels9SwmETHCwYUBSbisBTdbFvquTg7G
JvuV/g/I9eNUKpWQnMTHKu5ESXsWueBTo9j2RwkJwOoQd/Iawh71hgjrkuaWjWbUmAhzps1nwfpx
RB+/b3Pf1a7hUysxWy4QC9NvOfaa6Bji3rb1FzpUvHxbD7yc8rW0TfgGYx33exE7bQy60ivnpMtd
phxACOHJTJa4gkZB5J7KnY4T3kTzc5ELO0VmKJ9eduh7TIq8BuKzMffUSjQj0rHu29KBidC3j02K
tdJbsPy2Qhp1h1KfZtEo5kGvZZ5fKgzuPzt+1aXwesJyr4Ds8bRmJUdZAX6zekqgOdnlQIga/HeD
BUVcrhJSJiIp46llYlPgcqe7JXg+TQY4egTAWK/Pcm8+BI3YaElYkjR+igrja0syZxpJD8L94DgW
SHuGHZahfEZxsCx+nbayeaZ2JwGgO7so1aPGm6ngr9x/TxPEjbHk1zyhCtTp61hF+dhTBaQvDhId
fzvAfDFN2USd+w5CC/vPDXf3cZKz7wYr45nrK3h97kw/iPsdNYgOl3gdwMJ7wid8d6n8Sv1b6wRe
Zh1xR5DDpNAb8sOxXGf7mM6qBkuMksX2a352I0OkLMBjFH7P6VRzRd+8GtSY0Wlc7rxvAvzcsfCX
cMC5kvuDIP+CBJxXeohRfTp3g5aTZTWE2OXr1X5VmwrdXmOxJ1m/KBevUf7/KX37Boxg0wtWT7cT
NXzT40aVGouYvSIrVVodx/beqb9j38gX/JrpMlJTfn2B8ok4r9IBWirbDlkwY4y+DVFyBxySq14n
sg2zFDQNkLBIbEckrGVmDqnlGkhAhb/nBwfHYiEniV9oYrUeq60GwE0AgGW9tkoZza5eXb9Y5/i1
VVe2GN0FzYxwSnJakGd1Z7pdvJtGIUaktO1rZVg79YYADN9W9XPlCRLXhteTCrSfTi7kQksMW3Nc
TEdzggUGEzqtMPtQjPW1ucxk1Zv1PUYZfHAikweKbGbYaaFEDhZOdmvUNn3eHMsa9YoJKZvZ/gII
xCS5nMOY4FxP/Baru1Cb7BB+YPUny+kTzGmIi6cSkRuYinCeUF9FaeWuUIGCFNaN//n3Ehpr0/kK
RU310u/JHnyT7flcZM341STzFqGhNS7YPLBskQcF2TlUfPtXQyL1WCVfOgJvUdkhzzHeCC/3r/P3
dHREEswXZsbwww73d45CSOK9X5v82fhxyN2bQfpHsduR0LBaYwr6SJafnsKuxi1T5FeJSbVLJgBf
KrnkgABi81elfUpb+oy2lAB5rvdA4sM6XeGfDvrZj6cVIlXijYDAr8MSPvho/STKJsnUSskkmM13
dLjdRk5Ha9bxkI3PSlIFisIrxYo/i/fh/A0H0lXjSy0U9R3RmA/WMhHu2pZApiu41Yl/iRzaFkWW
Q7fjCGH0DPJl9I98Fc7Zx1ibA5XjT/K5v3SiM3kYbFZgkiTuNeu5JWYU3CIW7p4WbHio8RoLeaSw
EE9q6in/V4Wj1f2uSvNVw1T8OS/nNvXp03SReTvIb5epK9jLdPkvUZnhbm1TZRUPr5mwTebDs6j2
DoBZ26+Dz1BLmZQiW1mwgIuu38Yox1E84G+x2CFhqiua4t3TjKmBwVAskQw1uDRnfB36zL/Crhmh
ozGOnO3noYREpb4r4O9Sd+nddFAUbso3ubQP1rAtNRQseZYkj6zu56VlLCTt6+s8bKI94bUasOOq
2OaEDtH8wqVHaisQV3VORaFYinCPDk7mseqAIA0bxs1lo+SHuvmv3HJbQr7zGWTl8FUAkrlW0zFc
s+/iExLOepy483M+45VT3oJyeQvzE4Pufih/QMJGpOLeuaHbq+Icn/KGgGBXCSfhmpg/JeHX/nrD
olrf2MVH/KsIHS/AMoCZsd672E0L+Ll/y5yFpJZq5VreMKw4VMcHVEmdpCaZeFrEzInVfpNpE4Av
I1K0wh40cHnylQhD/Exa0aV7NHccmhGqKVa+B9PcsxPPQtVAvtqBbhNeUJ7KNB2sOngDQV0U+vQD
ss299BFVW6rn8fvP8g2mQI9H+GKcCiGuwFMlE4WI34nwy+ihzegwwVZaQBTb9FzMvu0A4rTDz5+3
Vixch1UacIcE6PUlAhv/OuiBdYw66FMkFYl2AMDc15r65CYqnXjV+FAz0ytM/92ADsUOE26yXcPr
ULSTV+7uaiZIRwoRDSfB8X6RF3Si2Sg2rVpoG01ooJngxjARlLyTR6FuoLpg8fMh66hc3rGJgFF4
h+q6yrP9UGEZ53YFQkaY4EBHOp/AL5brv2+Gf2hkWB9+I8/dFuvKQUjK/AQcJL0FxI3gKlpKmYPn
L/7AGZPTQ0kprjWvl0GczcvyUIAFznklVmTRENYODi0oRogu440qkshMN5hCotcDDJALK2mWVqVK
335DdY2LaoBDt/TQN04WDbRLiLLrCXV9gGIdkQGxNVIT3tONK3q5avxnmmHP7Ub1LbCVl+L13YyV
dFyCv0+1KYkNBkOCdjEiuhnPXTtsd0bmJoUA4gBEbxySD+anX+RL/bzefOK8dLeidw91lTGPDFXu
3Ui1ItKrIXH+idvD2RZuP5/5TQRowsasfsNxqKYUVNRpzLJdsskp7WlbUqCFCaYsPqMH5EEMF0B3
2mGuGyYVo5SAW170iZDoV1zXZD8CPFJQkZ6aNEnwt4TbGQ3c/OF8Z/lMKiY8F2fZVQT7CMbiE3q0
V19eDE8sJOZKeiQGLKDdxRKtTPMuXAiREUZXo9sPDUwJPvkg0LFXCEKTnf6BErKjin0Xp1/u95tD
80EdOZjFrIYwMI8DOL30o7JUXTKPZZmfaD9BVluGsjMCicskRCVmVY8dLfmtn8Qs98PDK0niUWWx
D5845np1Q7B2mastSiHNGiDkmpH6RoC6R/8dYg1VrZkOtqKeQkakeaJIsM2gfbA+YXDCzQMa6/yN
95DF/h3sOw9MxPfGY0sZ4XoMY+gPiwhZ1OwkWhAdenPf9ZKLXaBa1WJdrfAP9SK+QysXPdywQdHW
gCsedX50Hqxg3wUu4aOaSmFVhMoxytXAMvINEiGU9C/PgWhOmR1uazK+UY2j1kwboW0DgnEbWLwG
31Ox7JzpLNC6hf9Ssl/nAgCZnizQkqpRdKXyNHuDJH8Lggw8w+zg2RPnA+uuT1gkBbq1aaPxzlb3
myml9qFixFvpKAp5Y8sSp06L0zDtPrmrg88DvqA3rHCXvOqt+EBqDSLzlkNu6/bQkHeATDtl0BUl
rSt4D4CXyFcO/gDS/foNFT0bI3YHmUjrzwpZsMd4Lr9/LYZu1VbwOZVa34nyUPyqBHU5WDKb7fEV
iOEFRVA6EjuqsKyu9zzrM0ll/rwe0QPmj4WaB2EQHpQoZY5b7yemT1w3eal3nCrXUcewuHEpaAnT
Y0Fi+zzys28UM2DgWv0d3n8Mlc180W2D11czYCVfCOS0s+GIT3uMG+j0s1cTrVENF6QDOzGUdC8k
xhCb1yhN+8bW2N3u95GZvb+P2pPpM9O24FnfcW2XY7Y8pninqLfCBlj68gUFJDzppP7ZrMSrMeAM
e1DR/ghPOOBkQv1IiBQ1D+XlscjZzrrvn1H5vstkml0jcm3V/Lgzq4SH/zhtG/kbc1FQkxhehzeP
W7tSUq27IHCzHDFXYNtyTXEywFIdoc+lba/XMZjQQY8q8Mvfifs2OtpC/cXVo+0sF+BMjm34UoI/
95QIHD474nL6OaUNQOLUk1AixTA0TTRJeyneeYXYuyFO0Asg7sVvK3xTZNwg0g/IKO6SECAktsxd
ldZ5ffz9eKWhd9tLP5TbnuA0qnkKNZP0+QWuLt3K3wYmYfRKyGFDeYK2riWFHV/vssa9dLaVtQGY
gokVd0Dfs03Xjxv4pSu4TaPgp56hmvzRPzeAGJDrBa6sK7FPzP1I/AzHhbTRFov5GCPzZxFevp2z
0nRdDZff57QRUht+2jZ+iC+aj99cMcwLKg432i8xSTyBU4MYoljD8eNzy6m+AH+g3Vfi1k+0MIoW
42mD81c17gvr4gLOKpydiXMF0auEXcRE6pszo/FmVCMOyekBgdLTQrFwZkgmQIKtFQv87eg6RPTk
Wh9pHYISXBQEo6NcLQz05Bu1PLm2tyXkelWYX+8kq+zcS61WDEd7F8FAsgdYN5Y63ei1JUIzXVL0
Kyfl2DSyMh4Og3CHE6Vfmifjt3fG4QUXPp7g6DqFpFTMedL1UNclFeMZrXP37j8KmR67igcHox67
FuT4IjNdRwUXSD05YyViTjR2ygN9FcARPgsq6NMjSLa19n4oX2DozcoFZXvcw8mDQTHLL1SIY+cp
s0amgAI6I2zBvM3SKOFVxPxXYfg3LAIeule8YEU+rpWt8Yp3DTN26rlIwGR8OrhiPbXf3ZD3q1bk
PiUeubumm5g3nOOPExEMQijWOtyg5UBEGocAqsLT0Dc/zq7vwdnVfvQ7GfyJL/ucWC5a8lSB2alK
iRLGhVoOt7MMcmrDkLDr64d+bjWyyNEWXYsB4rVWZXVHLIaWqxRq4wV4qF28P/N9r7mE2Wnc7Mrw
E57FOI6QP6ukDCcdLqCSqDIJmEqqi9hBEQ5TRMHFBVwWCmBopIq1MR4qvvwoEUAeVaNC1IN+tQoM
knYw+Cdkr21DHLwJI6Ea9tAa2s0fnPFfI0oyeZzs65MpYakEX+WVwtQZQhruvGMrcOsi+6bFOR/9
8ZsENrx9UyeRVxqJcjmWdQaVN/w84MI0Ri1F06xc8Bx8CWjMZM0OdD8wjHymfj12oO2dnIM+A5AM
90OQciCBGObYvlXwwVj0mjuWZnU47/JYt6y1DNaZRxDnRv0BqS2GnapgGklpVWa2foWF8eWrMYE8
mHu2VX6jCDyE1CKyXTHDAAJsuKvNtmszU5XNxShLw90UusYpHxLlzWfIvhJi80EF391LJG9HD9pI
fNTyUajW0Mk6uDf4ZrbiEp6y7jJogOegYf97z4Xp0taa3Aa6eMCn4m7hV42BH8+mFXW0blVpVndN
fTnz2MPmLuW5O/vY3BiOlBeYhyRfD47pDo32DVrsW/+k87NL/0H3PFXgcinXsryLRKxZhxmasWn8
5SvcjIILjdZZ32WZdSGI0gTk3SMEty3gdxBckjpwsOXdAx2JWNk9x1JOicw3Bjf+5Npn8vjJ4jyB
FNd7DQmJQEjpC3gCBwpG4RCwPSN90H1OWzSV0W1atwg/PtPH1GS26bGC2TYo8kKVLXAdFnd2PB3D
G+0nUxp6Z8tq9p1zcej3xNBMJiPTZBpsz+cam7OB1/1NvAL7ftTbNoTnmdCPA0YhX0FuZFJe77Fo
kv/RV7jrbBMxTUf2hvPz9Yqy9q+IHSG5seqzW9FMO6yozbTksViqMNdOCEw/+1PUl4SJpbbK6Ine
R5J95faH64DxirNhj4MIViKEneQOnlAxceZodzAHEhpYklkvXRmkXbY5eIvy4+OLWTLuOWxBh9Il
0vQ1QbzrIbXFq2BrMPaQxdqPB9SLiSU20Lwc9RIoNOv8nfpnurDBrqvu2Ap9MABq65PL4Pt+XOMF
iXyuyAE/lud4RCL7K+v1WsNwTdtZvtRzRegbKex0olQbMhnjtbMuR3v9OQv8PyZmSyLdV2R9bwmD
DyfGAWzNV9Sx87ZPZbNoLYe+rnH9+fw151qhUH4MY9/Zmw4l/HXnYMiWIWqkL1ZbYRBIjZha6+aJ
p3lhJdO+8IuymdOwvuDAhQDmD8nW8ZXgkdVs1RF8WdXA6y/jSmk8L9Q4MdZ0ymclBIAqNQ9tIPaa
It8umwjtpeulUy53/6b9VurK5Ag4V88hsfkhjsL1ikOjh4FopX63SED5rxxre3sHjUAIK9xrBszR
kSGuIfy3Bzs2R5+lTyENOx8wqONyQgvGJDoW/hE15lsSnx9pCA0Z0p054xIuAy/GrAMHi+YFTdLb
MsNW07Pa+dTF/qd4fqws6lUKALA/mkWfJn9Y1YX7sYbYvgyvkaELJRWrk90B4wuMh1/rXndqVuxx
UtUqTBb00bLgd23lopdJWHVPGTG0Tr2Z/737BsyNLTXP0ATPAvSrO1f5XeY0ytpFXMMZSoDEJiy4
PmmdarsOQP8yix92//Rsnp8rRtYufaE6eOa8Y7vt0Iw84q8Z+bTgIl9quDCzCuIUQrvPtmahiKCb
mU4Szrlr158CcGslh9gsxXdY5zdwOSMam7TZJypARxfkMUC1v+m1zzFMXqFhTR9q/pl5kh/uLtSy
BrogYnDsUHeKXx+ooAf12y2vxnJlyd0gKR/Yc22v0Ecnpph3UL4/uEKZ8M81i3HbgV1WdvpYdqhP
NtvaUrHn7uJvhdHPBM3XBlNuqf0ntUEpD3CZaJW/7uJMjH31JH6uSAI3MOrKZnh1tTePYZ4B79hz
+Er4AuXmb+JNXwXYuh0yFiyiC7TYOuYvCN41fcheRP/TRdAV/0ASPBVP7O82N6yQK0bqixIgvXp+
xa+qNFkmwwb33QqYCOv9+u+okh6gV8Ai2khAnwuQVoGzKq37xqpbAdlYUdSbl/49pk8827QRzU6J
66j6YdYIJr1twMCYz0A+VoWkNZw2x/fkm7wLdqGo0dAevZpl/SkWk6pxrcEGL6ni7INxN7xrrTXB
fxuSbKWWT3uNXTSQodmWooq5aO0U+SL78CE59WlEZ+pUsb9i1KN1+x46a1zkyHMIQDuXWK4FunB+
UPDxWHseZc4fkHlWtK+T1t81zGR3CYxLerSbKYJ7IDqutep+tqZtOUby4gZou9P5INmqy3xb+CC9
bFbVXPSqdpCXpWrDFVpqISwPuvcXpJ0+lcp7JKcYD/M40uq4cvjcoC4P/ZIjjE2esc4WtxdpI+9l
MlzgZWgoRrObFPvGhdv9h2+SISAmXxX+nohPUGoSriHiRpKHfSvxD9Fj44KkJSTHZIJsOPygHYq5
lHwJX1QBxSN05YGEdkf5UHqCIZHBYlAiBAac6gHnpG+SOR/te9ChjgsMjKiQDXpo4k81Xc5kRNjM
qapVEkaGYwgepqMcGMoU5ZLeErp88SLr40vKI1c4zHtO2FQdPauQztX2/eBr1cnUZNh3h1wmsPsa
YwiS1vhc+3OOJStTh8zoTbZpIUNZi1txTJ+6CuH9ImOPBbIJpz2Q+LFtg8GhTyk8VYaM40eNX7da
rIIWqHHM17X6fw8g3PBRVdXz+Rn1MHxUW1UTQDqcZ4aXMz7SqYppdtraS+L0lDIGXkqkSv5RVZON
gZkVgiSKQbUZh1/jK+bIueTLJA5suuhPyWxu5EFnyBgZiDHB1ydf03roY6pnj6zhDcQtd1yAU7E5
Ti3FWwJuVXnRL9oAtsoRSyR3nEc/i3JJI9nQv6941scLlzkGjcc6gDM/Dna5LdekwdZ/8uduNgAl
7FppXu2aN+KowzNUY68tpEWlKFjdCcT3AtxUbcas63PZnxUlwuAqWRoI2OCsbQ915s9RlLi83v5Z
fnzEC7/g+6v8GpzmrVvaPymPw+sITMvC4evAqAT3p9c6pu8GAY6E1WrOB4KE2Sz3zilUuXK3dSAe
dufrc+pHy6B5uIE7aawIAkTiYp79qabe9r9iIIIMzhTgkZRA565aGcp15xQgBmVDytE3oZRUZ04N
fEVhgtUp3OEBBnHYGtCKRqG8bjgXypX6XVT45g7EJo8f60ANMeDbt810L/ubAn03uugB+m+rk9ts
PCyqd5loc10PY3zYHf0n5FM3q6Gf+bvoQB7UCJy5qsA0vbzVG9l21gNK975SrHiet5c1e4wodcDF
roP8dvIFGcoGIcdyguTiyCV6k+WhILKcmUtepWtDXLN9K8FvOM02726Mst9tiKF3Fe7nydg6K2vc
PDll0n1ijVpYkWAw7npJUV4XDka21zb8CYGPouCcv2gCVHUQV3oJqD8KhJB8/c047Q8x2AcNfVHk
Iw/HYUiwNvc+9aY9R2Wlk5caJgqvn3os0I+XN8LxzqcEtPGzDjdL/llL6Mm6KxftdCKpcyxAco7l
ADv2+fcAZ7ohcjLbZSZ1mFsXvdaqcGMQFvzllTm3ChORjMmyD1LvH/mvIzHQlb/0NKR87mM/MUoG
/JubPy28wtZ6aI3js+u8QB5O2vKZ9gIu39NyA6WbiiZnEX+1yIfhuPNMeJy0yp74bdI/5EH+yZ79
TbgpkTnqmQn5nynfYPF0mlureFbDfQsCbUOXQjV022Do9dxx2Esy8D1fFtDnEhWodd+o49iygAHH
tjPZvMOdXmVqCt97ltGXaEuyppcv7Jafxf4PxTGFOv4cHszirZnsT2lEgBbaC+lfJfrGTWVz3l8I
ocXPDwDNGKLExCZ6Nv2ZsdCSEOWwuMH+I6cniYAFC0sIJ+LcJ+WcoIBdI3ctniX1v+JDwhoMMI1I
4L0ITFv2AUqCEJF3KJOLYkDp6Hwxt3LUx3W4QUH3dmUlBmGgaXWtz1euZlFu05M0shra/OE8ZeVa
a25dvJINecoFlpjBj9m+ZgiGKSGU1DvT44uWAkvZaw3kmO0NGwxkh690XgLyoMVFRiUDhmdyB5Mw
FjLOrmz8I1MfAcOyYwD3sIEYzCHXVSKtPTPgnicR1POFNMy9S/VJsG1k5RO2S6vRJulgyb+Gl9VD
2G7IwmAVIRZ+iSlDB57mMjAGynixjGyqjdFFbzfutlu4TJBncl2+RGaq8evTQ6mmuN+FnAJj3qV7
TrfbJrPj+qxCBdpGyVDrfd7sDOlVIoIuNxUyn0mhJorLYvTKfVikSsmiH1klVcBGQZv2R0rWCC/y
ebt5nuLqrOfxJJ1ohh6fPNzC0HpyevChFXqAG8+POi1XqzKOEgA/iZTAuW4pz2p2Yh3/eaNS7xub
0vEpkrWBKeLvqm6I9W49lxfMd3J0BpILFjky8r1tQIgQS1B7cH7acpldJSSgrqPRNiCtFOFozgf5
koMulzGf0V8JIP2agNbqyrhzz380CCZGwWEmtUIdBC0aqrI2zQvJOPE7kN1nvayjDVL3As90SsHf
njcj77hsI7gGILVVJjRFaiUuBTTFuz4Wa1a/4DosZOR1OqnpbezIBXW1op6J2eAdSo0IHnHE49SW
WQ8DRrxJ47IxC0ixyFQe+W5LULzS+HQ1E62YkGxp1t+ol02Iv1mFywlSdtlqoqi7//0qMHZb4Spp
/7iAq9EpGWEKMZmpjozbd7hv/0YQOoKfsRKdpNuv705ZF0dP3qRRbZ8jZxs3qpR9gtvjPoCzx3yK
dHy+KxD3SnRjkIcrUzGhOyYniKGMcwLsUwLv5KP/IS9i08181XsDdoXh/bMf03WR8ceUbsb2LnfZ
tgYDQlppncGopt25+Fwa4G+xJFMXwGNrf1fsYaaImE70GA8ptjhkIZJjM83FBApauYqKmdwYU3Hr
HpOpSHekFIkLFOv50Qve3/puloa1zdvT9BvaFdzjotlsfGdfkxwEE9+cIpOrns3uUur0QmGfF9++
8C6yizDeagmGqbWy+HwxWF+BnxCi2Air/CGX8wqArbyD/uordTLdy6Of4nGttsCKHUcs1no4B1Oo
BCLvg/uKMkyJYT5umnjPKkVlPDSsAxgj2rQMMCB9/wm6AKxl6r4qCXuC85HAq9hBVFluTLgCfBCI
tjBQPnuDRq0k8QpqrwNcgojwBQDL9uq537erxBxtpW3XNfLPpIfkDe8BXyVL7+aEFYM0NW6K09Aw
t5W0jmGoUF4yLsDyKS4YeDSIgdvG7NqeVssVJ0azDxse85T29cJ0S03naooNUmcmeHqX9eKQVtP3
CxjezeXvIZaSaXnxIy3khokBiHDWugiBFAhGaEUXg0yASZjfRg9CtveiIGXpRSezzRcDvm0lYE0I
sRthcLHSGaZn+YcNhzcua8mcJFgxGUhIu3+pNluhrr2SsKkxKZP9IViBIwfiS1A7eUicG5wBUs96
nJfSl4UmtSMsSy//NBhSY9cYSCHu5J8AeKMEJ84n5Izc1ug/CS7laTry7On7uWwhMFskAxoEo+FT
1D8suSxcCXfhk/t1kZvPcLt0x9R8L+9m7PALJCqEMDBHsIBWSuvp8UPH6RYDeXDKjggz5ZZV79WB
n2P9kp5+2KNJ8OHzZHqS/PpWC0pdgkOaCAxsvvwyBPK9paRJPPV1fBkdL+aVNHdkavqCiaqvoRp6
JW8PvK/vNa8wK5Q7QyKpbrUQLoYTmupqz2L7pHR1ZEvImdCPa7VbCGRe8XRiXR66tXNmFNwgZ229
xtggn2TOUT2NcsYXb+N3jpoy9XRT1NytJtUE+kwQhriDWtSkV5P71h+UnN/Rgwv5pvSZQONzik9O
jpbv7JhUSrxIPTqii1sVBSKoWTNd5poWKsRVva7XWGMxRctmVeyWxaD4GrCPJRIBKg0t4codJxj3
5I0rDBQFQBDkh5tNj5UUo7gJeJWLiKyogar3fniTCzIpnZpr3+trUT0mQrV12MmVy2utUqtmeyfb
YYLvhVfaLgPwK+Xie/U51MuOgGixDlQe/5WYhD8JmlelalWLcbU/IbgKlCYuyBYNPj4ixweEySAA
A4OL8L716ZVi2S4P/StcmqgYUH+RHFnpMQANDRpXSl17tvYodgsGZjXADSM9C3W+Z7MorMLbExF6
6oNzf930fHO4iDHgJ+qSIPZ3ltYUHNYwjPg243v7F8hqaafYTARk19LkdTsuZ2HvwoTmdPIGzlr0
/8/rEvZPbBuyuD5v05PDL9N6l4undibiMJoLufXpsSrZPwEyrmoTNc8BJTdhr4YmR8YiaZp6zbOV
R/2AsN2e9jaX6FUcibcelmigxwYqMp+GfsmPdG17j8aUzi5AfD6aADUPU90AO32g0Qy3E3l9zjN8
GU+tqqDigQ7CeaKg7RqcF4h2qBcWksZRCsl01PN5gjNus4TLku2Sk/V2+Pj4UdQfpxHfAW0D3kdF
3CeZPt3eE99tJNne9+sdAjLQqpcrjDJucOHTkmj5jZjCFfXt1ol5doJzinnqN/FttR2Enh1GUlAT
+ZEc0QIJtRUK18YMETbaV8rEPkQY6JGtsD4ezdg0KWUvhz9it3DgZW/IRpfZVAm1C7e+T0qjzyfz
Wk5QhcyjO8JaQvpNlFvtL/oO4gjdYzGnBrjdmI6778ksaQaAtCxlbl9Z+D2ZspLF9f1bzfG4ydiT
PVfCFhzrd/82IcZRQyonH1TqMGkdyeXdyrpi9Uw0WeB3KSUUcSmKtN01M1CDMfo4OSeCVZJOzLuZ
IYSRxiv7s12JrsW/xJaq/Ovfo/vVkjVoyRmjGeFqmdzFwrkaIIZbbNLU31VeJ13LIEQt6jAIPWRI
uETClwMxayO5VIz6lfBri/oQqiUAtlrPPXv5amI/zWYWhxPDTc8eamjIUfiUaUWpQaRl0qwYb2UZ
UhpAFBu+VfA9QNlPe4/vGTuK3Mi8Nnc+nGpOKnu/p/100MfSD0PFUM0sXKgTkIP0z5jwrR6c/fum
DXcwyCkO/LlBlS1kO9tUPchTQSO7Swpy3MNjSAm0R0orkNorKGQdcuWxDS/z14mjKkT+E8LEWE1U
vuwzmIP1gQVKkxUFjkW8GiZNpeHqVIiqS8j6svA8fzwth6d9y0/YkkFEBb5zdIxzJNEK5EiA4kr+
h54Ll1pB3RiXeYtoA8kcVCqqPBowzrkyx+yYpLZLPydJYQkjLhiLIRe5XahuOypzB0T/Tyvgc2kl
sAYvCSP1cc3hBiyPw7oWYBJZyNnS8uWNBmFEnN6L2ufeNmwdnXQiqDAi0HMMxzKY32Cbimb1I5WO
VDO280o7ykNKHiaLp517YFAsZkbUj6DUmfTLxUoRlAKdSqxlhf3hlPVahrkfbF3/xGCEI2BHjH1+
PbiCt43tmoxdxlus/IlTap+FZW1Ezgppuv0LhmT7y8oF7A91lFLVfWVjV/xpYZvyl0QZrykCqFXz
nCgUordlqJpIrkrVCe/7cNAvvjWwpZv0nTJq9Ze8Y3/FZ8e8V82aoEoqBSpq0XHKRQgq1G6MfdmD
m2EZQ7fsZQUX/Jnptl+FR4wY6eHhrjE3ZD3GVUiypN7QNS2u4YWiCYaZN4dZtd3AMz7ISQAbgRNL
W/POvZlsVd22/fMMasmCsPJuOjFXlq7WDR1Agx2ZGIzFkcIG28d4xqih8JWsg8Z+B5hou70I0Dgi
C446/l/Lzy6SvrLqrtGaichm4kC4WmcBQDm4yZNHz7XVkK/ZkTzVDFLyGBYjN3uuOhVOmtw7xv5a
qs8zhL9LYWUi1c0Uitodd7aAfLhV9i2LbU5+dgbQ81BLNHm3oXz/CHggzAayjjYjyPLPrbdb65GY
79Yq0b1DkSl1/qY131jVlAYLJyBYAAHfXr+eUFJp8yDdJJAmFRatk+tzVPxtfBVp11mDSv/uh/7p
dlUiorQXvzh3QYBA8rRbmxr1AW+/ss6Sag3FRixD5PPT/Yn/ZQMX7Pg6CAn3J91l8ImaGBEu400s
4UgsIkNbaRW15GtG0O/uS1oJSBybHdjXkXsIrb+w7ORjManTbaALlVnh5OvY+GiSwDutcriL1Qs0
L/xFi4+4YpQ2Ac7JUYuf4Ccu27xOFSjg4oJLTuipUgycGV1qYZ7vLzhtxSpU4tZ6MM1NLaYS1Fdw
57p+h5z+kIO+PMp3fhYIqfb5BlhZ5RUemJ4kSgzxSylOJG8Wqppx3nkIoKpwUjEgAOG8ZTjEoEJk
GDeOM75tBnysgcsDMnQ43DDeEdCb3N3IExLcWF/0osEzysx7Anu/1myhBM/8pWUTr/kvwHH22bid
VS9t5TWCIglHH31Yzedcfwha7Z74ipHVl0K9uKWthLSTM2XRT+DX8OyH8yBfERvfyX7uShkE3/fG
yqO2Sks/wXrQyP+5Ftm7WV/ZW9OMgXKBM+n4YkdKAQIayCw7k9d3l1pMo0Lf1C4iYshvvNeUPv4u
LF52cpCDHG/FmrGK4w9Ad0gu7PstamazBA7/7z/2KzLEjoeTS5TuzArCYGJTmczFMkXoHaVwQW56
O6+g26TRHa7Ztzfwy3z4ybkMp1yS2hEndCMATX+RMj5LeEO6fClbMfqs376EfCaw5PedEevNDfCn
kgqsAwoX1ONgWCQStCMMjD7S1l/jOC0OTzXV6O7usAeRojSLaPw2oC/IFJnKMt/svTVszQRsYw6l
NW3V7y7/J0nES2smRkhKzHZC9MX67RixIjJmZUxAcAW+ktrXRKD+SuJ8j63jJZz/tP1AzrekJyXe
HFUR+xcWZzuZOPVN8AMvtiA0+Rz/Hwv8iB0Ecvjeum1sqhZPh+3KPpRHkM208ZC3m/YFCByLCkdT
l+8rj7RsfwECPthNSkK+UsC2JBzgURQwdIu/b+g+g1E104xbypHGiOTdqw1iZ0G/CE/qM6oYatXm
/vk1w0Y+krWuMyAwllouDh583oChHbXok7A1aczeAJ+FtXohx1p8wgPn9Es6eeqAnPxjrBkoFsaB
c720l4ipJzB4XykfPjUjVRlcmvxtvJ6QvSQfC6OwmZZoaHyncZcbdb44zuK//MIpUYeWlbacUEhi
cIcM0nDq32eqgE9mw2oqXKgz7E2+oWJj0qM8/FmtzYvCidkLJUr6MszVgwXTx/6KbH6U7UtJTUNy
2trmejq+WK2jdXVFeSkQiGQn3WAiyZI5m8mMzT/ht3r9XQFXvtUS6BQvr/B8MTGyPI9R5Ono4GqD
2ZFtuUOiJMEyuxnrXeknZtLM6tz/5cJ9wxz539IH8q0aIMAGkJ8E8Q2+ed96V5R24MH2kIRnAnUd
J9Rh95AZmuSWa7WTVF/qDXdqM3LuM/HvA4G8FNGEy/g6rvbmOb9ixcmhtEPekAYHB1PuHIs0557G
WBosDU+dyPxKoxXNbbu9cbIt9fpw9tpfIwaT/akJqo65Ecn6YcUPRu2dq6TOz9BG8bNz8Atc4SY5
si730f4KFzqc0NOxSMBojP0jHV+Ad4s8uijy+3DreP7tiMstJK+an+wzZiRlCDnEzC20WlVKPZSH
yUjaRdbK3ue046ES8CvhUr0aSYzAx0AJq6qwgDvVa8hel48T5C17b8ZrIhw4XJvzfpirQesZCXh5
YI0tDEOSzMQ1LX3a66OpuwLagPjwyMwADzfQvG+/41ECrZ/tbBqq9R8eS3fZb0DDkvvMpx0aZ6pc
0ImTpDcaT5FVfYQk8EDI2Hq/avTvTqK/k8VWohggV4JKFsAPVXQpqoVf5ao0DXd3pMUJj6SKUb5V
CYA3IvByYIhW/B0WHsNScesjOwOEX8fqjhSlavon5Hu8x0yzxjbI1Zg1RTpAT6o+KgB4u6M8NaBr
EVOfIKBRbQu54c7GW0a7nlNa9iYik1OFL5GD3IFNFLlekCqLq3sz/VeQT7F2p6JJc/wgYSzUq3sZ
9OMM6sokegHRSO5mdch9g8Sg5tgc0L06RUVcmoLAp/aZOCCL46XbKNUvqrAeAKITWpH43PpdmcLF
9fiieHXcx8yTfRrQ1RcR7MGBgeu+etKhJkMRJ8OxFpYxDhJxxLa41sbKlbIPLl6lAdwtLXkO4MSq
sonKpWuNtUaosWGTyzC5bNX3dFLLEOxAbLe53JXejF28Sdz5XeYc0ATduSlzXOIBkmRL4K1LE7+6
St0+2p3/93QZIzE/49B7atbXcQ0SULqL6EGRRyXktXeaJ7q1vdCgM6wgaLgGlLsoIYlblzpbJVg1
39awI52sQ5+NgGH179UjwoSZHzlOImr8qXmQjlJnepq8fGvyxlbzMCdKVbd37p0zzX2dzF/MjxF3
qGGPJLjHuX8rU5dbXGBgtaCzmMGip9H9CM/w4NITIzQGauOvHQp2UMqa5hQQUgeV57uGQ+XdcmP5
vGGaRa7+WJFExjrYb0ECmXmahxhtxVPeMmcvcUqScFT867x69JMwrmjjZmdWdT9OvAHc3lYs9UJn
ARLVAhMgB1FRCElzZGWu/AMq7yb7oc6xKGKw/3Einl0dXzy83alFTDR4wg6rXD9xvVziM8B4cg8Y
29JIh0s1vvjXTTDO0Kvc/1V+CD4kmtIYK5xjZCWwtYIv+vNsU4MFVgL1OdDigj9w+PYP+d1TQZqw
PC90dPzaBR0UhbCdSX2JX8Y6YdzID1sNlsk/mqKGvxNCzwjyZYtHYgVa/0F1z+zAJFxo6LTp4ChH
wbyOANre8asT84VjBiWFwO2WqUdNPtRwckLi6Zchp+sGfUb9cb5wpHHy3qPagRVnI07wFBwDn/E0
xjSOFZh5TqZohR6X/WmJejY0bahqKp5H9LIcCRyS46peR/49fPXfiAOsgHmh6Ei1m37fR3WOAGen
M6sTLtHA6T4P+MPLWBbPVJjH3/d7PjNMXUDdoGmkKz0DqmBUgRRVnEtadMblCEy9iiphq85X+Ydw
563ta9XzlVen+EjaosM3QdaVXQo0s/37WLTvt7l9BxADAWtPwqs7NCXMj7/sn5wAC89p+QECARkW
/kOoVhdQ/qUwfvDujq3ZpfymoQ6eJEolWOYZlcYtEJsHBBPyLicn1GK67Sl3DTUz7LOEf0w4WgDj
wWb5Fxru8eFmwmrP/wJ1CmXgnMUarI41NNbFc1zbQYn5xTCaF9fjobzCp7kYeTMA4+ONrfbwF4rj
IZd7t4mzTxCyb7aV3FEsJ0OWInJPxRmpiBdRh8M3Rn+ThOYYECpFcUQIbuMjj8ECssHkQt6Z35Oc
WPrVUOPpLDUXaYErGSefy/DYZsy+QCFnzxG+CmuJpqAUudeeNm2BOkgEoY+DwgLFYiLcDSVQxOt7
nbCgyuv7fe8OCMgZSSNGG/bJYoiE8QZ36+1+sKrugQ7VdeFK/PSmS5fv0/51khqioOHsaXoDDB5V
tmQ6BbXablmJUElMkgAICtvksjvPNA1El/2mE/VtD+kAtpkKObFt/GAxQGOCl6ubqklbPosi4Fpu
nGClMPcdDGY3ECL85Ce6kcgfLJYP9E1bKRmq6C57fJaIonNjQGPbu19JwX2XwP6d3JuxEFN+jVq2
ZsFPJYIW0/cAhWeZX+m8GXnBmGmwEvUnrf+CQKfOOD9JA0mn2b8xcIT8EyFw+tSi9uVUs5R4KDPr
7ejoq7nX7/H9rtRtw4deO8U5MY641UyUJoAajMKBiO1/HCuW9wRAKBkS2Jk9bJy2j8RPKFTy0OEJ
3wFSqgnaYKccSGS8xNCOEa2bnXmDCeb4A8FJKmbQ/NtI5NfG40QixKg2KoN7Vmkw2N2XhibbjvTo
SaQROGFp9JIhmKHfOXxLrgx0XimrGZk3jblR6lT6LA78wrmSZldE85gQVc5nCb9w4WuKOrQvxfuF
mpqeFWqXGzOwZLvhlmmRzz7TFRD3xmMd+L9lI0uisc65DYxLwWMnfAu02ejDeLp0vXK4gBJCamLK
m2PqqOHrP1z997KfmJs2c6u7t2Z5OdQBU36cdgaWeGbCXISHB4EtWwSrt+Ooviv1boIsIOBu53kM
IRu8CbAsbQAeIZxhNU5K2w+btBEdw0/kD/vnXV2Xb4pbp3lkTY7OIMZzSMTsP+pC3iDyKMYg0Tre
uZLN5QSFLLuyFK8Woj7xvVVbjMJU3+QR6pGlxoUBkpEQySN5nyR9/kPAWqRj9BbJJfDJNZnIq7GS
rTI8IQmiSfUT08Z95mISnYeIOXOSjaV9vOKVpluseyGLqvckMyU0MNnekVQw8Q4X0IBX7AwK1Me1
ffEnSf8AX5guWyGoxUJBNYaUSeD9FSl7ckGCLrR95gYFNUv3SeOZT44PPhMJxsfbPccQPudQ90uL
Jjx4ABTJ11IK+tSk6wZRB3Ckv3WvVMM18fNA22DzMmAj8oe5XMQhpcv17hegsAdDxxl6XumUXBaI
T/tg26NZ8/wqJ87lqC0JneqZFCLjCEZ01tnO/7yYDDI/9lk5vUEbM00GvF5HG8la9sdTCk1jhD4T
OA01lEsGplYlK822zwzNV6+BGHggobtE/U3GaBJco9miIt7buItQosLOqiAZzhTIq4zSG223MsIO
PM9SoiNH/smEF+PmVAtmbiHhpuA3Y7WUudANl/DO4iWdQQjDfANdcfD9v8j5d3DktEXJrCAWkUl3
0kfBM3NqAT/OSV2joLjury4SauxdIFtwQ7s3c2gekYq5kmiMNRfTzXQPx3EONQrOfSVKKZXeT++y
06YZBG7uikUvy87uqUgA1cSGTpSLhVWXofgr/XxuqwTkwSdBMMzQSP9iSWD9l7mTEWsjBI8EJYlo
aUogZbFZe3zDsz+xg/Ue5dYO5Js6ZWdiDlp5bnFMdlsfoBkhAfGnMZqvE2Sl6du9tLBcJfS8MXG4
ouCMHhZVYqPwM9aKfs8rW8qdiaW6gu47Lhn1LBV4Nc2kUfzYVBvkKxD5dPr7aI7Jilc3uRDI5qiv
iGLiLC042dnrTKQA0SJiXT8aSoi6yKsCIHa63eAjKoqImMMiCIVjfrarUsBk5TUGdQ+SUTL9VaL0
NAuIfQCcB50SkxlXCBLyYdPU0ilqQK4/WWJ2Wqt2potL8EEoeqtb01Ih2zyjWpWS3XDhTutCBiOw
gnKIE8zW5r3aovzx0eu+pEm25JxYMQRUCttuXlYq4Hj+KcUym0Id45O421yYLsha2TfjgMKAVURB
MaTc0hfjMDYbLYYrlUDp8/ml/6k/v090Sbdt0wXRIvCc/Yfe3o/0Gb9a97P3zZ4AmYIGYmYG52m8
kHw9148Ulc+I4X7zCr1o5Fj1ZKmUUdlIPI2lYpV5ayMv5v7vr9MXGVHNUj03WzWXja+8bzeBYHUr
vwl3z53cmsWRlTZbLrC4GVEN82hcDSnO1rVcqB1wIRw7gXpE6XViPu3O3vRQuS2qDxsyv11TYMli
b9hdfJb1gWwOAwl3YAX7fGqP1eOC872iOjDArip1bNpHn6QMECAM1r2xnv9D9rLkdMtDdfffQKd3
02qUvL0cWiB+ImYOPZ2NxjFe0wVf6a5+OI/7E4R7X4xJMUVE7+41jdDTu4vqgiPh8WKR3zjPhunf
uvMND0jlTL5Yb+56Y6aQYkWufW6jPAVOeH/yIi2a+XsYBSg35u+x1GkhYvDcdwdv3TelHLSFmPNs
cONhC5MbwMiDF6SGPjd8HGgf71YgX2PTuN47mq0AZQASTe5PetLxd2FfpfJ6eZQkL8F2Kf3m1F0d
quDyIfRnlJuW0cZ6Yr2ph48zQgzmaiqNyWqemIS4fD2ePe2y5N5zDgf3Jw5oA+ETJLkrxdz5I2fm
elZw6seIFbebgxRiXckakjAFpyPc1fDL5GtnMvXzPL6s5r9r5d+03CwI5Ee9WialGcXnswD4Oa8t
n90yAL9jivXcLjwQyYAu6/I84s6QBI9mK5W/IZZWSziyhyuY+zsddhuBw81jYcDW13l09uFQK7oG
OFfuWXY1lo5nJRxI1VR8OmM+wcmjA3LNa3fOzsDqDdKAnhSCvGq6evKLt2AadTETi+4bb4J4XdHk
i8Ib8kTVb1qUUMaEZdl5FvduTUNW7/4rFQSDdiY+m0AYjEZsG0sOm+S14bS+7ZnD0oRLtN6Z+ajU
JsL23sbr5RxmLzGrvjpkswKvhkIrqkRRLRtq74FxbH6OK1UIj2S5ADTw4S+Er8wA8sgsHkNFSKxD
RwbCXzmn6np16oStHdSUUMiiHuCXIy62wIdX7trox+FqZ5tBYyrejwGmcW3v6uwHajZx3Db4y4i+
CSGHzHWOf3SL3lkaX6IQDfRg9xzP28jQLj0xXMhwhfI+AzrbJUIMpYP4J9Pj9VkLb2buv3mu50bX
NeBfvxBlLuVXOFvwqmf52jPmx1WLQinKufasnDbQIwRBQ9KRk1KXSPx/dlzxpElSqjGE+T3XHxgM
GNfcF/Narsukw3tjvc+jrFYvHdQzAR7m/hNMFhJVE9WTIb6GoMWKh6vkdgyFfN6Nf/FRk0+l9Hox
N9a1yMeR2odI0MqezclGNhZKV4XFdef2lpRP1QJ4Yn59KGwoTPDmd8lO0kQqxKpXbnQfuMLm/Stm
KMpkH1qNW3fvAGLcm2IECzBDsd+9leSR4vHgNGkGmR3zlE3+fVkvvPUpCav8ukmtKpswN+4oa7+X
x6AInwN9fDaMIRbLk9l6hxVP7oU2iJNdFEbwKfmcvdqZiDsieoWj+I5j402rCC9Vgn/hC7PaTKDa
oHRxqZeOeWt0XTXFMFVmwPTkIYStEQ/ieQOao7EyV2JqI8i3Kt1buh6QgxmTc7LERqCfCmLCcDyM
SANrxWkS0jZhiwcwx6bdj1QkTdC/HbKZ44bQKfCFxrc+CTAQLKthu1xBVMcDgJCCJ6+SoHxlcYtk
QMwazm0iDgGWJeRGXDI5ukwvaZ4kMECQEMIQZK5BBXVrna2JtWRZ3u8Vs/i/g87SJdXobB4F2vFF
eqpGftKjsXxZfmilFrvZDmV7w+kYblJVojRDwdpqoBs6rDh9skZAfazDiV/MfFfmJoG5P+hN2K2g
QViYM0Zf8mVZjx0Hcb2R4nRPNG0orBkckdPKCIKZBrOEaRRWna3hQCt3qYHCDpZrKn29OSMQfCfG
5bTn37/MyBIzjh28TQoKUUqpZezzyd0uuN97jgICFsJnhhlBNxxCOHTYCIgnkhkg1BJD6JtF46x0
Dvt2AbBKrTX6Nahb9dpXK2/iJ+MirXSLqH1CTR1FM2FPnVTN34Mxiy5HaSTQH1qX00wNUiBoGzTI
vwffAUTtQvos05YxfP3Vq/N+CVXtk1v3woTPRpK7ZAlGDhpTAVDXoTngc5ukXUgeQYY0k3QC3a44
Jvb1w+ZhBC/ThAlu9PbzlwpXKrATkMyinUSpT1vE7OBs+HbCa5/y51g6XndAsCP71XfdPs3+h5NF
yA0OOgZSWwbLnhE+XL+JtjwIFwcgtWGG5VEcSs5tlczDuHHjKpUhNkCqC336HfP8d09C6qOKPzhR
W5jyn0aKEn+lGIqfH8oQHiUvs+HWM9gESf4W0a7wa3YtiuATOEo8K+RY3Aqp6m4arbmMTZQR/m62
l6iQw/53xHOZnXZKdva5+jhB+3jmym9To1+HVCeZ4J49g+66Fu14IGzVNAv0F6OkQrwOZcffljST
B32hxwQymSDAmcIzit8XZbXdxTNCRpR9cpKqosAzb0jQKOQXG4zI8JuUhK7kN7dMKyRgmiqGyGAn
iBTZ0vuFQM4T2V98cO8lZHGRLs2rAu03tMU/OeEPupXN8z6sDl0OB1AfgxT1HHAy5+yJHxueoLkb
xrE06ccXdVYub5JXYJH5t0wudQky5fk3bZWXDmUBQ6AUNNJPA6pw46SIkkvdV+y3LbN2bZy9My08
fmPqLEvSmvE+n4MsjaCVOjfzV/JEWzfcrzugItoOEqVbUqyrrX8syw49hk1E1YWQKI/LNOjDZzeY
37IG237RZ7M92aTAIBDeZpnAicrLRODi+zxc7HssbCR/eaSCDV9BXah5IcBlFQ9mvh+WJqB81jXP
MGwFkltiZdT1djmuIZ3Vo0Peouq6JdKYPRxwagtFtIHE2huKrMz3qr0at7tFX/LHrqTu9a/NeZ8V
IW4mOOgyWAxCCapPG6mi1w4xVdbxWaDM09yZVhvAOL3mpyEeQeRuuln1sh9VbyUGTbkCXeHpvBRp
zQpKeXKyq4AYjgclNiQSo2PZSHDrPyLkLCfs/BOorq/KwveBdnDAkJUMzkCm2PyPm2beBavnfLER
BsrTXqM3/NUOu2awFzUZr4a2IIPVOjb1cOFxFj2spILZC7SX3lgmYb9PtNtFy4YBhbCltO5P8GZ8
KNu4yAVhj60Pp1rHSQpbC1clIgOcvuM5ud8xwAfcVp596O4n/pGgrFIfpmQ19UHEiqnUw8ngoumR
YT+7eGqC7P/nisOVbd+8T+fevDzTByS3YJ5a72V6x4FNfzypBj3t2vS/64RHo36WLsvh8ncW6Ph6
+x4lbc0kzdypllaXdWoDGQmp5QT2h1Rf8FCbTbO2JNI3HCnZvS6o945LJ7RCYLrRHaxNA5CucE1A
ykGD9nIKb3tezl0mKp1RwIwvqgAsChcHY07kcdEVuac6jxgD4AmL0NQ6tbvru1jR45qolAR2kOvF
V55NIrSH2GVonUmNGYmM+EamgIyE0eqkpKKk85mlBxreIUMuOI9qclwOphkr5TKe223DT/Q5qXhj
oMsG6fdrRK6EDr6X0UyH3KrIwxUHArgYO/7DsDV1b5/bONUzu7rLLdxWfGBIBoooPqEkdKlqnYeb
wkotKRi9AjAQQrD7EBGmTrQWioRTS+dXTkPQDeEInVGkQrgGdUgPfhA0Nlp9YGY0Ik05ChqRbO96
8ZdDNDnPPGJde23dMJpEyuNxGrNN6cd3IRidB0jYUOZ6XOPyD6ZU3BuWPeLlqflpMSoQBQMPp/Qz
TIZatRLsrlDXw1KAMJS77TpRqJSqcnA/+eZaUp/aedF+WOWhN6gS7fkf7Plgqam3pZjGjsCrWPrW
F4jUcrs3fQS6SJz80742rwZgdqq7m6CRgyZ1RT1WIKAMkrZUdBLhIPqunvjZoqszdooz05c9D1Ui
z8lT/+k/ZqzIatIDt1LDkD9rKCLkEkquIsyYvhGCfMJ/gePLedusT3G/Ra/jr6kC0meqC4l/j4jr
fhFGOMfueEE+7I3WVg6Nr733XLyi+831fphi1vl7Y39vu8DPVAryWKjjmDsh0ntQ956py/rMgkcj
9bHzRy6nOpyCnTb9wjGDIPQYslY7L8sF6jtid2HmYM+xAEPjsKU+ZS2FFIZ2YgV0ornDjESW1Xsy
/eCStfNJ94zt6LKzmBi9oO5xsuG/aCgeb2t8bpd2AxbzUcaukcRZZJnGbwmAapo89KOfKonCmmpK
FIo9+otj46xWQX3hi5ncliedKt6qyhgAcfLUg5LWXFLRKrWTQOZrvRbP0n/5PLAwQ2rH1Z1hSnh1
2xID0XtofjQChmSvnYfe/Ram2rDN0zgSWIwtOoOFANU02cfAfj8vTvz5et5IFZbnScnVXbq9YlhF
7y/rd2xHS69COnXk3P0g1+5oV1JkCdgfhhYl1Ul3VzIu91+Rs5RmxHJo5UgCURU7uJ4VlOriL6nA
HjuWoYjPi2DRb8rLz9ljONe7sf5HZGBq3O8qTfooyWALdKekBBnY5IgfHDAPJBuYircI3jHkjU4u
HoF0B+470wrdZClMbuSfKOGP6pPI/+hAkcwB6Inu3+YfsEe0vpx/7V87UsqI9vu0XIteYXYY8bX+
1BvbMYOxztoVrytUwLUau2KTmfMn+zDMnExDYOTt+DHqzP70BLjpTz3gYqOe2wbx1zH9p3Ko11FK
Wi+SLw5yFaA7B9xz9JvpX1XhGC4UmJZ5ALErNgAvCCRoWrOlrwwGTRzCQKTSvpgtGaDV3I8wq06N
WXeGevjPxkMHqtltV2lwof4O83vWb5QzijzSs/bSIH7/OExgKQM7E8eyjqP1Cqc0v2dzJYHsORuo
GzwUDS96adYUVS8bJabstSzODm7guVijr7dBZ4nSIFF0Bv8kuJLMb8syhcvvuhGPtHst+DLg9oHt
0dvAj5JBQ6u9NWxfUGZYtmtQgTXO7lUgAsNkKU9/zv2hn4zNIw7KuUcsdtW6z40TAacavJfMiP9/
F17PPuNLwoI84pD7d8A1DPOpTq/XRAvxSwMI3ediUosz3Bw2QjmDJvcc8shhFQNYl7M2pwwSwxT+
Ngz714ufsZFZfnXw5bY9v6jCXroJ4jwA6RHLAERSd7pNveRNo3NB+ZsyNcyZC5C/wyX+vOU4ijsw
EnzYIDATbGXI2IWOVdqiM5JosaWmvr7LXk+NVJTrtQgrkH2CVbmovUpF+bd+Z1Yv7P6GrhSHmzA+
u2i3BbTUpg8Zj+NegOmi2p+IU2u0lz/ar7+Kla5Vu66dBLPR2jHPMl7Q1QXzEl5MlHwx9vfAXRlD
Xe7SbhuXmpPqqx6pcFgPoYqGI4YxX1g5H5a3LVE1bQOBC0UgHE6Zk9G7WEWJaxQG8ABvJ217VMmT
BB+3vQsevCuNEIHNcMdCstJmmnUUmRRZecSdos07mevv8ChJ6T8xCTx/PkTZIEtm3zjomK6IC9WE
Hz88/cp02tmdOJ1ITWLNM820Mkb1o1VufzFPBcZCh0lGGRcvAL9YbgYPktxGorf9sB1zrIQpM7BF
/7eTHUKh9BA2Bf8e5RsCjs9c+Tf8Nwzb047CK7+UZiizgIFnEvfLCvoeQFlNWOqaR2VZVcMlOguc
Q7tOZ0UA4xyEg9iv14RBrI9cZZIc97zbBBWf6oMKIyE5aELSUxXZbLlgvBek1kgkOcItu3/RywNx
Jde+sjxWZT3/WVucJkoCs9XA9u0Sg7dM94eUgAbbbL9xY2YogA1KgkiSpTfnWblFNjxROWvScbBc
zx2dmN1PFnHYQdsDiq6ENMKTnxvPzs58t6ZRjHTELhX2HSatY2NPG/9wigxw9qb+w42jVLmlz0IA
Sp1Ilp7gxnpeWV+JtfFIFiV2MwUkAtAK5PmJMbP9OAbVTykF9nJzZsvQ9DhIa055f8rIoNgtjeQq
qjigzTlC65gEckzVxD5tIdllkIaXcPTEEYsoE3yoF+4fROQN8qEL6WGOsNozF0GvGqzdQhCQe/pZ
Lw7mpSVF1HLogib8kgXWz1LA52LbWfLACMx26B/Te7blWKNfyFWSsgSADWoNihVg52Xmz0HsYXYj
QPgjHeUC8QkzX4EISQMZGyAfBOwIG10Sz3lG0x4j/x0j3tk+2krEIUXWUoz2HKlHK22BK+ZRJXJp
8u3Hq25L9eltBITj79K90lz9FTDl7YqzEsPg5/IFs0ZUzen1oY1JjcL4N7ESXinhydBMU4bntYv0
9VmPfrYHpJeh42y5hwAqY+cGkLxf3bfVln4PWEqibhaaOOR1u+xrSuBlaJANaCJyyk9zdc35nVkx
P4rL0KV3Oid2ndZ2p+CsLBYWEIEt0Oc8meewt297BHbDxcf0zsE8Ms2fa/D8VCVdwqtTeLYPlouP
oapdgKxZzxBqWsibctHmFsPRzxzcZXSc9RvSUzVAV5EOXQ0P2Q7zJVEilDrAg74RKcdoLHkwFNIW
wU/ozANVNV9pue/pssd8niFe66i8okBEua1BfqTQZWVuSu4KWNf9VseNlTJVnE4C6JtRCB3Bzzsg
Avm7EmuxMJlNOQwk+SQLUkUie6kLAJCGtA8Qm1siZMr3psm/V82C+TS/9qIsGHEhGY/IC6FfiYM6
kV+yR/nGdkNgH9WT0Pta4iIFgrjiE4gJJUO4aXz6gJ/nTVYzG9NHT/Dew36JVF9sHwllhDw9Jvb9
EqDq/S4Mu0bgW6aGQqfwarO+cvbBJNOZPEQ8bYCCZm0cVKgFFgqmKLajbJ6c0qsWcKsOtuwnIiBD
yy1QLuuG/xywIhmBqTgM/+EV0fOqxfTE/WqO55DMEHFVS2peTARutsUGDdUqc2ab6d9JY3EeMM2J
1ZuLiYv3IaAhWGMB5Ku6Jib85zdmPjWVWQq1WLRmw16A4XgQbWlpa9V2nYOoOVwl1pTE+LfuCVNr
YLKxa+u7cvuux/BLtID8oORxBiVKVwMTH2tlrZB0TCsCiwgnotm1nVerJKKR1h1oGgzsh09Bho6m
RTnu/bguXuoiFJudZUWZhd8i9f4brWLc0VdTQSwCZAoeyrMescNFlSN2SNBsZULTLcYbbis73v87
k/mAGh30O/Ab7beZ/04vQPwE8l8zg8Zs4WGggLLgOoTJju+24CXtMIwI7w3aSgdw402VHtiVNdtA
FB/hAH0w7kTpYB6mYLcb0oeMxYNQpDMqfDSLhkvoppVb1uABN4KrhI1+tNkuOHlskz2cIv8/dPvv
S0yN59uI3a+8de61eZLaGVVkA3+xHHe5qsGUs2IWXEJI9Q+H/K9XBleNZ0Q3igQ+7E8Kdmvx1Wvm
ZHhGK7PBwJDSaQq4NZFfpCETXpD9AnV7UVAul25yHRxaN0WSCnBufYs0PJcDH6RMGPRh9JNvWpwK
AxGOFLF+0wcR8wfSY4JJWLuhRUPmyKno1eaFy17ncEpPkOYHyl624gu5VZwKFeQEYNhBkY4oNh18
NyUVMSlqFU2LWMGMqBYW/twpvSoYnviv1+QlaQKhyKOjt/7rm/3VWcG0iu6hHe+6jiJhVcgPrmMx
vqk7IjVuFxgX9E9n8x8kdZY1DzRW0+zJ/bp1dNFLrwhEaw122GLLV2/XlyffEIe5zQ3w0KUnlLNb
JVZDX3oEiCberXre1qRJrtyyTVcR7YuYqBdD0LefxVmJxHdARR9rk3ZgusGq7ObSaUIul1IuZMjP
l29K3z/gwLpUGUubrhX8B37W7jjOkt8Nao6rtRdJ7fXUJaKBeoiEFi0AoT4R/36JDUgn/3ZkolO2
e4MwlQxk4fxEFs43VmaAd27/iDOWrhU6wELkVeRmLremnmSiujFO4P8z2KmD8YhsVw1jbMmWrIus
vZ9D3aaiErDIqNNDR1QyDQ3UnjwNzOXPAAhEBJAQXgwVKYImECo2XaoCZb+XC1JiVFCB0eEDOIVK
KsAvaJe6qGt5fMk9SVGG5vCAYnsWfd2hY8IsCrzFeb7NsrAw87TpLpGIDhgSX3mkD0c/A/dzez6o
lSoQYsZ3Ps85RjVfB+yGaYkoj2Lri6hFbR8tR0u3Otd3YK9uzFCLL5kQ6A2DJncArq0B5eFe1Zgx
znvS1WTAweOSpA/96G7IWL5ILli64qwGzO0oq6S7dWzrBnub9SG5PjtFXFlnAoSupn5ErDf3X5Gt
Sj98pT09Vs+FSNxSCuXTpT1vmP55fetB2NVwYPmqQZHT7p2mEldL4ZU1ACc3/Cq9RypkApfs1USQ
Wobm+TygaG6yN369reKU9TwMRORa1dqelczzEq0hkBvaQ2lim7UKNngBCBU8r8obP2XesvJ/Iv6/
RyFw4e4i7Lg8iMW7jkfReHhRD+HPjbpjlZhEJmpT6sEKIJ9l11P69QameZ5TApOAuIBkfkFN46bM
lw+PYdJKnzksoXUDv0vdASIOgyyk4IOD9pRFslvW2Q60MKv1Rz483vPl0XUhuA7ou0e+npXh9Ba4
atUNoqzNSfBo73MmZJmp6ccUljTWjOUYG2kH67+19GwSWsJTJ+Es2TZ4U7ErdUlbkycthXkjJrYI
izyzB9/n3YUD0IWlddEJHmbTcK1Pp9np4iP0gYMPlymB0yHLO4s9SCT6xtVhworZNOQnrpZQgSLE
6yV1rlKzmeWkdBlqRiQ/FB6GB/G1ji7jWdwg7GBAa20NcVDJxQdw/VVCb6ftSpS4RAtFlZYvnHFf
kvIFbykvJr4nq9jlo2cBVCpv4y2NN5dhna8KAzQNYbjt1HJiSpTwB4BjW+fMvoEXcmgqppebSPQS
zF1tMvSRIq68eyq8XclkIu2lxbuPGb8Uz+CULivzNKUL8vyEVXLUmOlX+xPO7F3nVzEYJSY7oK7j
aZ4m5jvTARoRJT8L8mnOfsgnaxYewKL7QE8AWLC5zpLr8tOV9Or66iTW+LKvDXwPlVfkWNiVUhnq
8+LWF8QDaEEwPhBlzRJkUTmg5qs/1aGs93D6TRbEIeNYEmG88YB7dG2LFsScdSGq5sMPph1mnrgN
j+t4nZO7i9mtIzqGKgOYlavY5ustRYb/4rO15ST3947+ltYPPDExg7IEzF/oRGyyhFdTQRPlWRga
GokVtMSo5ks6Cl+l/Rky3KPCdLP1XXdUGnYX5u43TbkLOHTVmmDXHS6Ke/JFEXQEL/mLhIMNzJOi
CL0vVEwP8Va+yvbBvGMhPozk3pZ5LXVPb1YRkvViR5V2smnVP0XqLT7cHoqzCbe4Yai7t/5cTx+F
BGGh/pD0dR/KvINT+U86NLDOClmsKXfT+WCdH4Ebncmz0aA8FA4NvkeNgYFO8ZCMFQpC5MBL/kYe
B2y78yA6V1bolB2vbrognZUO/qf4oM0Fee4ofZqxEG7KeVz3dkps6W+I8z8A5ieSPkJOX5pvzS2k
3E7/rYlPXomH9eoTmdNZmCixacmw3ycOEMJsVWDA8gkiQnVkUMOuIJyySMYsA+SxlueAdwW9Oc3O
zN+XkuCnAX6x5xoC8zG6OiJ+DWX6QCcyJ6XV0MEzh/4PTioFwtvm8/DG+6nv1xTNwZkGcj/Q89V4
lSwJ8PNSQ5qEkNtkel2ZyKFpvMkCk1fUqsfUio8IEoy8FMfTX3fxiLHGz2NPlu+Lft8DCJBXMptA
pYQF9/fSsbMwVj0G2wk8LzLHoIgJjiR/e6Xfh/SZLhdIag5SQvJ7qOyTCi28cUWQu5NluA2l8Kf6
q9WgQLHiHmQftLUWvZk6rlxQuGvI/V4GIt4w0cUS80td06tveJrFlja2NNLvN+awHRUY+bXD5Yph
SNykvciDZZ6CIestTqcXQLt9dKac3ITp+0sODXvVNQpHTwOyqi2CpS7iCnOcnaMytbPkTvs6o3G7
Luia1wQ9cysG3i3lyYUOrz3bp2FIMQzgsiHeNmpHuPhPaJ6+vOh5UP+RneickGc0t9EZUoDJYaBi
AqH9m3ZTFLb6zMuvyZBReIDbI5Dr+DuRRAueU/lvU1rARuC3VvjTYK/iSjolhis9X4Br/sHZ/Z20
U8QDvLg3mOH+briMohw82pCFR729lf9+lUEE2goh0piFDQobvAOkww42d8WmdyKV2eJULxIt/viG
XK3rFSGdG2kFyzMD2XT15GsdC1IQc4TEIYDrWy2RVacTOdQh/bDIg/09Atr5DH7n+5ZGF+QxVFSR
0h/WDaDF+xliymQysRaj2bOIRKKkazrtB6/HDMqBEF9dAwooQfvWfM5Ub0mQB11Q3WVK1PoNsWlO
zxcXUeelkNY8QLEkrgi7agzhNfPOTWZLY94qbsN9xDMNVAwM7+NcXOGFJ0cMO4ndZQC4QrruQTuL
+HHpOTzb7pfNW26rYAWXUJyvbz8zAxqgAfVKXh0fTH25LaYbGXoaE751PWTqKoGJputTYSvtw3KI
QwOetwMLMK+jyIzBMVdSvu0qlqYHbTrMDuX5xayzPgS+mcsNHPM0+qPkiJURh4GtFiyPmZeXao3u
Me7AlrkT+jWR2S84VwZOcxFmAIoQ0gssXRAIE2o1n7oeK11MHen6pvlJkiDm0+wsGVJD5Wej9xfw
2v07PEo114191B1OmAcmRe9/bGIpzv1VkBnPN3v9OAjmWsyToKTd5p1WnVwPjx6CNv2xmcRjxWea
NE+go1PuWlUIHJpLgrljzEQS6qLVg8x39a6BHBlva+/p3nb4NLxc67BIUee8DIxSR7knLW7OEXzg
9hskDMZC9/NUMzXnBTv24y6BpbjMygY9KW9l05i0uh9IaKF4jwLhCX3DeLdHsVKHJDJTKSx9prsG
SuYxvf/9rZpUZ3OnXWDE2cVJqIxkYGro8QskjA8xNyOcYU9lTRfnJoQzmr4q4BtF9+M9Vepzdm0V
wl8C/gjG1GY9ml9NdqNcsGFAPKiW5xIeOeBvrSTcLa4eNCwUSLrlCmL9FSAmY+Bi0nhxBsb6BQHi
gD68UWrZIVD0ZselKAtYA9ZmXMP4qt22ZJmeopovFFilnJ/uJD8xm8gCp3G/3//wVZ/N3OnF5sW/
wM3Ko+imhA+G3ceeoO+hnnH/NHDAW+krFSf5mKrzioBrXwNttnvt3gLP8UoS5//501KN57+gMKDf
yS4IQY1FUBLFa1rnP91bK7c7PAuH0co/zHWJjCkKPbKoZa4RE7RLet+gzq4xiX1LkBFu9kmskw3E
GF8YkuYPKX91L6juE9Z6gNCxu9GhE3GeP0UBB17iC7uuDx/JySgFWiTP7+M4sjCDSkW5O3u86ytv
ViJkxHHD3WbHXsOvDd3t6ebuGkGtGHjDFJWQLfIMLm6LyvSEaQ6VK2uf6E+opmr0hblRG4+Fqr7h
kBAIGb6juROPQJ2Oy/y2vCEKKqIT49FpO/b/5BKYeSPWScGMrdrRg2PmK65/GTPVmQtNRnD2huaS
TKlwe8x89usLWvjUYMPjgopwYqpiclv4R/67zNml2WVkdLGs4ulhkdn4vedR7J0fz7feyatjYPnz
wxDkegh73vT1Czk6Kva7VCvrKmGQJcspf0lzB4GL9GCvaHXAknH5ritJr/eFWYvOr9orOwZwtnTM
6iUzUnqDflfB4xfJp+1EgnPZFb/DliY6ukKYDJ+PyXDHRgrVUZD8bFlt4blQytAKaxXzJG3vxvPN
bV0E+n4ltrq2BxPEDFANF4fORmsKy/hyRwn3hrs4mxyI8EcWNY8v98mNHnjAFacFg70YjtD7/D4l
Lt1C/z2+ZXXZDIfSr58pgnwzDHXTKdu6sbFQSUkHgCU1z2dOC+4wYYUklqpzetHgL+Yfbv880N/e
udxv9EWTq9TH9E+WjLoM7yHSwETQu5hwsDR6dCn1pwkFHXGxGKf5y9CX55o52IXUERupXlW2tfvf
qZ4VYCbD6FC0liOJlPGcKEBBeRyHsMEuQ92YDDCKLTwBRdhI0lq42M6ErCAzCrBD3RsLt/ZB+cdO
KoBNuaewhi4ZheIfaldbRbCU5iBJdI73hSO+83HrdvWl7EQ/7s4uIgTFowwpayKeObq8xsph4iX9
jEpvVocRfG0GiIpeJEc+NNXIif9Fct95Kv25t5pyPA+eKDxcSs1d1e3a1+R/0AR4EPhFSWKQe4+j
TNHzTY6JbMxGmqnrh9a/qqJD7BrWJuydCqK+KT1PYCpubJOOcrFfXeb4J6ADq1onIvFvY7Y6N0Vd
heH9ZDZ4auBYgG7GL67v2c9e6sRVPN6tTAHJ3pn3Fs+1UrHxK72yt0pVza17k8kyjCWN3MQktcI1
/AIRZ921RQQyuGjCLseTJEDcvPoyT31yD2eerwGULwweymlRlQmaxrQLiLytIXRYSzWvVRJLBNEm
5Ll5HqBUKaIiaMx/GXABoDCzBmeKjCFj/0Px1wyiO9DDTiXP1xnUgYKpI5dSFkufQnQu6jJr7HLk
K4p2R4bm97VnZSEp3u/ED+MBy3XxKMGsZk223qa4ofRLXU2RXBcbpkE6muxcdolETyVgb5ESpie3
RB0Ax3xYpcSMWYjovbc0QjcmGBl1KsxFN2nABELhGQ9QNQd3Dmm6m9GxPq7wT7tojQeTbD/rf0eJ
uC+PRXhL5NG6Pbx9olaIRRo0Ku/tgJuq+cA++ZKeomxc0IjdilLCjs4BhcbyoRbUTiKVOO9J38uu
i18GIr0mtOlQDTcV4hR0mC+QYUc1qIJO/kyiJ9BW6XLzEIPcaS3CTt8GRvtbUyCwAfmz2LSqKSIC
bHy3XBYOY2Nas2uT9Obe9zPnV01DMhD7RyKEAhPG6yBBfABIoWyceylb7W97CSM/DmC4XHpi3w85
I5fvMc17h4xWOrJOJ3eqghp2MYPJsz8Vny5dTjvvGW3v0zXIdIk60R/O82lGPsLgG7oawx2Slsbu
Oi3SjAv+v9vA/wAeOoZPkCamJLdxNYpMns41PQjLyEfgBhV/wD6wPKXJ59ZE7U1iGD74dUpPzB8K
jK51fQr0S7Z5NBq19snBonL2gIkHRsnjOvOdYPG8FMdoB+KGusXnf0UMf6UgGJwqoLiaWllBbAUf
gQkQrQArK+jlFms772bm3Ht6vtY2k8ESvkVWeCfSGWl4nEZTPWFl1SuiBoV7RyEIVFX1lNZouKYN
SplOctHRb3fqAKGd+DdilxTWm1zzQCPCks8JF6EMLItURRm6j7I6lE1vd5WdmYNvTQHBVa9U3TAX
F2Ltwq027GhHE2tojdXIeETzWosIoymW92mY0Fpf1vMH/xSGrYRCkmLBcfhzzUKjt1kddmKdY76W
ZOpjt0+vRtLKFpuM012hcKkbujqgSpElHis5iaXUAdE9C3a7WxAriVeBTYZk/UPO1NVMZX/WEulN
FmYbvMYxoqP6I9o2STql9LxAp5bI5laMQKSLZRKBiBgxGKqzQgQp31uNDekNlcAj4Ux++MZUXW7Y
fwIV8FOiOt7V7J05jak8wlJfijo3IHPM1oWbWZX1PG6f05qGxEky8U7C+oKDXJhTVbQCh4smHqu+
FIPuhlxsFxzLFoadP3RINL5rDd8FkAyYyOEyeFP/yq+jTfQyt6f2pJgPZ/9U1PtFP5pydpyLfr5Z
/vwHezUL5C1jh9g9lfBN1JyECCpW2QoWpQjq2pqWrOepBpP4cPQaiIzJUE26YISuI3vvxD5+FhHa
zrAcBhRWApuV8YKa0BqsnWscN06jT7PEyNjMBvEy7ZJ/pcFWxHaWSJU5skWNONNqP7JwqVR7/uB+
cnE/WtBRBxCBKiZokyjTS3wrvyExsoTFgfLHQ/c6j6me5G89budvwrZcyDt4WWSKgISuhPy+8gjl
kPkUw0ZPdGK1wPeBr47N6UYXQdAcbABfW0jUvKZmA4yaDsZSh0CwL4G/rgJp+e/WYxGakc3KvtnC
thxwhDY7VboxK47xWfp9JGGxeo6W3LhBiua74fX6Wp7blA8EQ/qGjTWCGK4dVqTmytzR+b/K+uHw
uc3fuVnXVBMJpFnq1f2z5zwngqeoIMV7rON8rmKZj9wRPuk49I44yHplQ0tSRHDCL/r39RBCOON1
9NjSu8wWgVUnk8rr+Tcgkxb/F7C+zdTzVchdVyV8lClogvmZe2GP3KEy3aDRQwD0bjpQBTE9FebS
8fai9wjA2WRR6qM6jmhW58MpPKv5eVcWkpYMULFAatw1Mf+kR9pttVmXo6yAVwXIiY8CsrKsNy57
O2ZMNmVq9I44ZdItjwH3pKD39G1wvBkPCnbPG4S/58S6lnZLzgTd58YpofeOHSTGRjQiwaBLy05/
8KGUZY0SDhuzM5KEbF38AJxJArz3I9/1jEw5iL+iX6O4XFh/wiih5O702nW9o6hZ5Spr5lrpaaxw
hZJa1RorrVwWHh5zksGg+Ygpw5aa5G3oPdgTBYD2MJK3btAEvPhoalnCi9xrHcfhC23+dWo4igB2
4vmeWLx0HH80iaxWv/EStGXzKJe3/91ftUnBZL1GUneJcYgcdrkIyrIeDY83L/CVf8+MWjXjGuLW
ZNYDeY8CdNT4p9RbMxdRJVd20TwV4HNMToMPSLVfvcnUP1vpEG8opydOkINJkSLLQ66rMDgFVASc
VBlRfZqxA1G72rA5FBAggS9PsxuVfsISFUW/lGVpez87MdTrgUi00SPzVNZkK+Z7068fwbLfWo+t
kJPcScyfFO5Uf/mw5t9sJmRcGL5xsptcCKHuczDm6kzcXJuHy0c8VuiuyH5AK9m4lyYVq0NzrLNI
sX3Kv/gKB7Cuq4qo/rQHfzBALqzCuwlTG737CtkYScR8xqk9FKFNPNEkIZv1mx6Q62tqhRCZxpj5
G9jxBmhfib7NXlpq+6n8AZRqkUkJo8rF2TVHE7N2XVJ84j4Xlmb/lJneRuVeS6YM3c34mj+n8YIX
0yWlC1GIp2TKChaeecpW+y0HvwM9O/Kcz+oRnvnyPBvIbyBBRpHu11pjUVy1M4q3BlmRMSZV3M0I
+yAp/4E6EoYxb9aGKQOejOiMPzSurN67JpWExosJSmWXbpkuOyx0goQ0gmfcotH8IhJtJl7KVjHz
nxYrR0VmF1VsjcHC29G2ob62BPgLjrzCtBAd6V6x0RHCqv9Db4vSJeQOuac4pi+dWPqJIqnFVdiS
jId45ls84H8O7/ftok8T7s2SLDsKxlsfxxY0QI6FpUNCY6vYS1hPwkq+1z4k8Q8knpO8z407aA/Z
FCYHAxyOL01Ras+U8wlOGxRNijXx8kCH5DUP1Q/GYF68wLi80O40h6sC8kilnG7d9DWAqzLz7c0H
nIKMix6CSvl7STNlPSxvYa5fDgj25O5P+fm2aU0yc9gj2Yofa4IPH35hv9rybiuhe4EocQauM9PN
RHaSAiKAvVSOdvH9zrSscL8POSpv5fKfxzihwRQuo+7e8u7uFR/zus5vwBtnMvxYhU9GUnkwu2lV
1t7sJLhQ8hb8unw2QCuHWFqrPf+edEjS+ETaO7KddV3aVrw4o1DdY3umex+7K+ovZzruipy7Y0IX
S7ZVQjNALP+EAvXTaqcJLfV1rP+ckhjsKHyvqHxUBymQTff92l9I1PtseKI77iNvbA7A7GZSm8vT
ujxEM7ABiuQTJUh0Im4C9fO5Rurltm3pvxeCIIWR/euo8tPIBkIse5NtgcFNxAk7DMIXDWh1XNeL
QPr6zFbWYZqOwaGOT1GQOo6+xac9UVg/9CAI3eBXAueUaZqtKvlwZZtSrZInxSaD5jxVaSYZbg4c
f1u+qXbXaMP4QTc5d+hLWt+yHMloo5HbH6My3ZKiTWv5V5Tp4DO8tI4who5IdvLLuDMoULX7Dr5P
xP0KvPm8eeKB4TbqGTVwA3YDmDBMktY8u5EZuN2dWe/NS6AXTysT/v+z0u7dkNy2dS6era65qkmx
A4Z8uHf7vTl/W9gKZY1YuLYzv7dI3wcyNopyqkq0d1gc071m44rkTuHc+U3Y4O5sCuOoLBq1hSTE
l+YLWQbyuQMvA0Xq74hTh8c4GAGjd/crkprq1xbx+1yNdl1mHj//N5Anj1mWVzCAlz8EKwOjHtut
/lEL3I0GS1w2n0c+BrBoEVZyX/JzlvyZkHkNy+9z8lMx+v1YoB1NRjjbt3WUFvjlo7BsV5WpTUyw
jzp/osxIF9j2Cs93nvd+exVq2KZxzJUgduVRxHJu0fgk7fG1r7AfGfkseG7iLM+EAFn0b/SV5/nb
Ek3InwwF8PineXTd02I/9xVY/Qow1REh5p+HbaYY8AR8Dgxq4Jz9vmB3KFFvZHvD9Y5Tq8CAM97l
yZgZIM5KMkC2qCKuYXHO1RemaK0CvV+ztPchRFM6BKdxNaVqIyPgpphjl86Q2Rexq3GUTtzDwkCj
rQSN3HZ2oAbpdh2hEUsKWHFp1ZdN87X4Yng87M/GOOe4lilEvqF6l+MDkVlyVbpFv4wtQ4dzo9ng
6NeLY4NJzq/h4j5nw/dxRM8KEMSKbRQ8iwOXFTB8sMNpp/ywZqnF9ix+OgCls29tnMN6Pzq3iJ2Z
/VDlBXCXhiUtJINTAMeZ6W6XtK5W8VXVrXPbzu41GTRHU74/iYZffkZqmyLH0Nj7d8AUOFlykQfy
XYz7XwYrVz4iZHQOpR259nYl+OdkII8Ev9DvMEMalhxenHYl7FxHI+rdSvGKUg3N5miU0bkmSFp5
AMtTnERTzCDbZuoy6jPN7X6G+BfkzK0RbkGpmvjJcNrqAfsxTjNxBnffOSCl7gTsdT+pk9bPLY0p
o+bkVCYdxQIhPIUm7Itne2VfT+JuWx7ZYrmMaECgTDR3kaEYti0kh2ho7PzjLc/vAJTFn31MgQMK
Hcl4aHmZfPOa8z+1JZPKfuwQws86GEMlRo5aAtG9teDtF9Tm0b2GBYy99tXFfHPYr3XBnZgg2X6b
ZCbra3tEtbKx7GOBlvFRnO+liECsw1zDNJXZQH+ZqtGzPm0GyIZq2Hh3vBXtpeO/7g2tEKG41qwZ
SMz3k9eJpJBZcH0RKVUnJRCrh5tJ/6qrR4wW/llBemWPeHyRSn5pzsG2O+h8qiyvjqVMrqu6z45D
oFRAp8Yw2VtLY7iJ/DiENWbgOgp1j4OeDoD/yOqk2zAxXmjXFkpnRM5uuXMEypMubVS/q4MaT3nG
CESiLmoQx23P2nfRh6WxnwsIowsc54+KPBYQbypROX81B+DmIXfvz+46JWweXkCOkLVdGtrryEX4
fy6OrqxmEaNo6AO3YpFtvnJjduW8I8yBtMg5oG5SwyEgoCkAhqFjnMvoGrVq1aX0w8eAmU2QHWAH
fCkJBHU2hLRKmPXx9Wj2cNDjhdmexBAaMmm0bEZmwp/NiGhaPJhobB6djLZVKGyJwFl3oyD0wvnB
UGQXOObuolqP83k7cJkvbI7PO1zWaurJP29/G8VLiPekYbJjrTBlBO1DHp66RjoUYqSrQjZel+4M
9pjc9SWE+Y7mIwrkn+rrrtvg8v0VuV42jmnSnk8XB9hcwM0kiYBYoiK+ymIUtJjnyQc6RknUPjZg
vgQp3nWuyX8wxSfYKMAkJyOFlVmSr8yYjYyxr2jNQc28liiy9BLvErWLKCmWweErMHgaKKewMw3w
XJCS0QqhOCMFoNXyEugS73lx4QR3ZjghwwNB3XoJzt8RRJqCT2qxQQungWG+hX0TMgu1/MJCea+m
HdC+8n/5PQ+UFqiHm8SbYdkRu3QH89isuMthxHE7reBXf0V+YvTCa+YT7LjsemAWD0ZKiR8zmXP+
p3SOeOy/EKSCUZOZHfcNPR7pnPFd0ihHvlT1018yf648x+EjMG9r6Ad3di12yIjvphCZrCWMls2p
VTEmcdqnaJAmFzj+7Z0N0E9h13J+feOHw6Tkjlpp7Y+KimuPbKtjH2CfehyQA8pUpwNJkA+w5tKd
LK21XSCfdE8cHcwDbtbEAyxrwrRC1Ib1oMdNgwqKgJyONRpLrKkdWsUio/WfYXVEQ4hkSIwj3FMq
YMiJQjAxKBhfZQGIw5BaASfv1AuQ50oOv8Uh3OFzcuCZjNssyXdMhSl/bcB8IBiq4uIZU9Gm/LoY
2CtGjE/hFj8uFViAWMe4TPFA+gg+0mW4r8ZdgoIKmuEpCM8DGYb3bJEpil+3QAYBCC9n3fkrxsz1
YP3To1JtzjV5IVRDMTBd9JEIM/kjIX/pT/odpoQNHG3K74zVj4HCWWtyLMFewCK5Cf1I3+Cvpicy
YAvvVdj454ie/cInKaKbUPRMwZvNiQ8+16GVqCk7QKwrF/XIDeAZoyaY/RlFzvDKLOgrSpRJiYoC
e1LDrV7ZlpjqvuoGkgBch8cIYkg93MaoUzh1KHtC6mSWMJT0PeOfCa5WkOckbsJbsOoPkrkvyc2M
wALXSpGng+aUGXsqbzb6j2yZARkO88jagGQtHdZjPkmNGxCcMvT7bn6yC4o57fTSFfROyJtY7l91
HUiVTLUiOqn/Gd24ehwyMsrrLlgVbQRhQ6kgt1UX0FNYGX4DAMdp4p1zkfoQkKQ1v+vvJguwcNmy
GDfTAz1g6e5W7acsElIlntd7Wg/TKIWbqwyj1d6Ao4IDHeI8jwUbd9FneTD4HJAl6GuFFKpK4Ll7
4JC/h5FjFgYrqNHak2Zm/mggMaZ3EYPaV2e1pilQYupld3PQISx7UZFBZHUBlu9Lgqu1g+Q5TxPr
rP+78YHvFyUSTb63nYsV6Iy3beao7CUNh/dF5EjvWyF55wqCmFiZMHBHEb2pqQgn+EwRRSylDf/6
012B7giQdju3lsaE59sIWbzmCK+uBzXWYIwhGMHxWAzN7JNgFFBXqY9NffxDrdlKiptGY+5aTQ6f
YB1f29lC52k0gSxPYKNJ81pMyjNiL/unB5Qdr5uUwZfLiYvTSeuxNNO8+vCArak1R1ZNJKAzWAW9
jMiRQhqMSma+yyDhgmUbO4hbTrXXNhhoAFGRBKqvubWSUKu6zLrv2auyl4lU722e6cDR3pOTXLRj
MvY02+MI8hMIyf0ta0ctH++SghMmYvyTqvaoixu0/YBrvw+3JD8ggGEr8qS/jkBLST46rMpoBQJO
yP8mmlMzJonhmCSapPy8wLhXN2FufzT0F5zO8R1S1quN1Sq7/EJjcfAI9ODPecT+SvzF6VONymzk
S/RHy9zzpoZpzxQQ8DcUzXaknXl9/Hhg2fIMlHNJr0u//hR7yQiuplDiCwcqdRI8MdkMFEB7dp+h
5IN2C8Qlym4aKNskIXal22iXVJzFgqy/FDFsrAvC9cZ2IdE/N7ysKdPYX5EJzWkViFyJmzKVgfGO
qatxlf3jYRCvB0UkG4e6AL6tYw8yLqXZ3FQiMsPpNpRp56nmtJDuym4/K5GRAq/JbPUZDO2xhQIt
ncUqZsWpFzP0msCthZL2zX50XXfVINioOVWPVtTZEHmBI3bUFebqk7IET7QH9DlSJ+Ukx7ynZmDU
8FzUZl0EP6VOMntiTpLx7iuZNtADbABhCTXid3tur2hCfgCHN5cg5sLrIAKfDwFpsM8nYSYC2HA7
LjdQhUFbTkvvJH1T6OlPO59qJ0s8FxwS3WXFvwt+o1v0HDEWkSdcCHuDjisz3wVECLjyBMJ+5uFc
u3wRA6IX1zbnXR33LM1jOxaW7JChZAwxHZKM5dpE/59QFSaMA5+5YYKC3m1+Nu8KkoP1nALA9YHY
FtbCHXnCfObo/XfonNlpPSPAhHPpXuHS1LyocKo6A1wzVgyho7PWqELTOgkQpbe7fhtssqheEMcV
bVKhFKRK3H93Y35KWY7kPh1aGLQXlbhmQa6CaP3+iNgamEn2FeOZwGx6mxFyoWIIWKqwd69Owk3j
T7Zd9WmNMrEVV890ThnDpkWWOynXL1iLgpT9hQtQGpya7p4xFhfx8UjwSQHJ4jPZUe1me4zKGRfZ
wCkedMJIiQTllj0yk9ehp32uTtwl4GMmlBRijxliN+zTkZ/alenLDHUngn0FeKZ5p7aGEPaRmLaA
fZKyTJVSuK+iUj/nd0FLqkVBlQDiCM0deF9ZY1/whtyM2Qeac3aA30BpXfnK8qsA4V5Gd/pYRsSN
hq0dR6wZrExKdVSV9+yTDZy9KfqVL7VX01Kq4YRKn7q5MXY/YLOgl89EAFnXeycxx8P66G478nox
sZL+xMlGr183Flhni968vAkuLvOsJ34JnwdzTE2KIlgvGFny98ui6aw4YMsx0t8Br/Mm6L3iFvR+
s/xZ04pgNDx9QgL+SrRLoKdy8M+ALIT6iwBvjTlQb4wMt+T5q0mwgyI5aTK6QRS0BTIC8qcx3GPP
QklvI3dstbPFTYfEyR21qABku+y+Xla37CjB+u7olU+jKcs+og7ebxRqn2dSy5+hQZFJpV+LfLl9
4Fma2Aadl8/W78gTR2+/P9DYn56iQ2NwVOIu4LJbpm6XaJ11pC7v1czhmPUBpPQPYnZkKB07QNgM
KMqY1LlYxo5+YS6n6TcKZYAF0u3THVHFhy+M5rfxrfLyQBTV7cyQujpYqkIo8xdz5KdS1S6ehuCH
wXFewJJTj2gHynNwmBYvJ+IDyE5GdJKPPEJx229HYDcqgT0cSFkCxKq+tK/96uhCFoubgYCdGai/
gUFwA1Oe/bGVRNzVkRAUdp3aZtxmeiRqzTqkpl/6E+cQGVbePwitRQdQHa/zSLEmgICbsRkHnZ70
P3/S05iTAYe5GX2yCid+GKZVatW9XUZAaHLFGu+1VVl6WWBacQrXIZaVBPXTcy/7DuWlNZ8LMx/F
o2vK4uxesFww8JxI801Oq6aOAReNaU043N1cwF/GFDQtOWi40RrYqKfRRMfpfif+LQ/svYTihxn+
/vG76Wdog3PHV5qTiArYNGjTIeOeQJD1vzETdtggSpQrvKj510L1IwgQ+S3ZHc67yLuiGq+J8Pgf
oGw4drjxxGkLXQdkquyNMANJirYKOv6TUo0U96Muq+hFFLWR0Y8C/kEFRdgB4OoGJZXfybC44pXC
hB051U8NTMA2u1E143rmqWlmbZE98S0Kg7ylGVSXU+7TItz/wjL1IPU2oLY99DmZJeTO3vSgNPVx
VoO1h89mFjoIcDZ88rIvNO1bZrCq5y2xmZ2chAw4cVw+DSv74MLHN5yQy8uzW0pRaX746t2UlmrF
pxJty6LgxiodyC4VJVdI0XHUBB9bneNjheI4vP5e9Iq+UOdUZlyHyPf9pOghCJarw5INSMCNIIm4
wpt6BUBEV0Nym0LLgx1B27s90WPTV6/PXSro6bVf8DNDHIWn9nkTbdqC6sCdL4z80ZtzEcrZvQYR
9fgXk3INBUYn922LHdN4M/vOCAOefq8fV9EDCyW9eYHyiMUUjP8i0ljxv8b82gSusI0HzuQqzIIz
zsmneL8LHrZYrLDb3TD6h8duqlZzDawDUbsLNejy5drEU5yqpYNjiZIxjn7m87oJVFRhcRMmijPJ
HmuyJ+ZJ5TpniIEfMZEBE/k12e/qDEDK4qCHhHtA/lFJkUiCO6v+AzGvV4cmWOVwAHmfqPgNyb3j
zfhFADdmgrXTmq98RM5X0yBmyvAfTp9uqvXP4tFe532GyesSdgxWKTDiD2WLlVb2gf6Z8hYAL7Uj
ofl7EsMVS1K3ComuKNkFy2H5cSE/xHOeKfTMEXnIbV4Z5/gUrkFHyOV1OIbaJNbBmzEcpTDpoGhd
i26iX/ab6nI/p9t21fGC+rKdU5glJ7+Ai/HrqS3t+JtgXVps1K31TKwhHzmniHV1wfNMKmADpKim
g2OxJD+wT5FtlDDGB5itUoiJcEhvTLodZB3hHWFsEiAbrQeqgpSKy+RRgdkX2fNVb+xNDkrm/9tD
NyvC8GjTBO7/kCOtTD8RkTOJ0WXsMqyPv0tnf8lXkYhXaOhsXcWBFqFxMRnZGUxVO7zjLmY6zh3z
jggwbTIcUdPXyPUxuiCX8Ff0GCFOaaP76ajSt+4JYEjqwlOPpxjAgYMxwzlh9Rh2I+HbkzKXVHDi
13dTuz4DTjQqSs7AjRTaMiCwXADEJLI3CGKSf/mZoIMql3LG8ABOg6jOVJjQpZRi+WTkCae8Roft
zrr6A/467qZ8tVfP3XakqDWnm9jMaBC3q5eLBVacc8StO55xmvY3XRKlQ6Vr/xo6W8hoSVSGC2tM
jtCJRYeU53kGOpUsV4RyBPK7t55pMcG0FOlgaWAkYa39gXILifyfba+OWBCkEjD77JS2kic9k6UA
Aer+9gxeF+leo3bvbYd05Kg9ixH7NC6qndfKBVCzZh+SEAPprd8N9j6SUZD9KgAmsPCACQYri+Ln
V0B+jsq5KPvNRqFJxpdQrNu9iGwBX+IqnG3wEXVRfgHmEKeWUlXuIh5BxL2n0jFCbjkMz7467R+R
wXnqE3n/K0mQ+fVfoi3YMuB9DES/KjGLwt80QV9wxSVc651EwmdEgQUyEbQVTfYleYGR1TkGzGvB
DfsNwnn0z1S5Dg4+5+9zQVrO1FFcsvYqdlZi9mvLbedmijjFnGJkFiKoqbLwg1rnakJ43n11Etxq
Ir28PWo6IdSBiFMD28b3dZ+EOKxgNR9erDjzCF0Yt9fTxQPgqmB3JPG+Xk6nn+RixIB583/o5epx
99Os9zjjCbgU81BAcTalMC2NNG6guOZ93zI/jnlTV+dz9UjHZF6seRo3xEUqPqyRtVpdL9No3VPL
g+/tNic50QUZlwUeB4KU7rO4Z84Rc6d2ZijwefEpQlg432FkRzyflZ810k1Ml734wh+vm6NhvGMA
gldWmHOB7TsDNyvJpdBAGnOQxZLszCgbV1zDs2k86n8OsJv53sXffFU8aTZGWf2YNK4vM4Qdza4t
TTUG/+61vGzNVjRwXiFYC6yjm48v0XWkZMHxAbuXSilM3R6fFY54rBjAuGCqzBcpelbO7ZYbsZoO
y/k16+jA6SK/ZdlkJ/L5tdUDgA4SJz7wMwHZp801HYnaCw297SNQusKm6SFk75O+eWgkgvTy0s4x
TSw9qz4mEVtHp36sJ6T14sCZpbrNvpPOvnsJen26+EA5OePriPNXmPs1dxnzcrJbEP3ykTu4AgCW
t7OnAqImeCtshImUlD+B4MG5FbCEniL0Qn2lM0ea1b+DsmqNJ23HWV/qjgsKvMVDFQpBVLxZ02aC
KgL11/S6cXHKfZAZn9sUkMqDRWTfOBDq617fhJSbXXb5fdizSB71GU+u3IhK5mENioJSL3v6Y3kZ
ARjPz4TMuZPwRZwfDrbJ/KH9e+NxneG+o5kF96FgVYhfTx2ZSaPFKe9/f3iAlV9r7pNHxBlUWJh2
NF/KwNaonAx8fhMrK2cAEJHHuRQEC56XwsAk38lMAUK5pUbCJRXKnBKVXSfBkLJ+NMe+3R0z+EA2
IKYI5Yrzfse0EtY3/Kc1ic8oW0cMuOhDUXcfGcKMpSfUgBpLlYmLyBzjgVe3G4ttH2aavN+B5Kmi
m2tP4h6NaLKWovR4bYrOup6mRRl/jb6P4N0SAYY4W0Iwg3DEBy1vdK1TOsw4fJR3YdFXAHUZ7yuO
mFJew5PFf7ojfxR2KcqnIEyWTPFgUoIRKdkx6tT75Vl6FIsMNhhC9B3HDnOXLmztI92TQisVIGax
GvpCh1wgHeWDW2NBVp/8UpilGsZAxXpUjx39d/WuRI+lfEFAK5y3OlhcTMMHSF1HGG0jtHbNI1ZD
sUCcrXcFOX0pK8biChhCH7R/mzq4ZYIS3WuuvdQiVOJa5ldXo+L3RQ6ufP3+j4Whppfnko2Jj/Xw
RVSBOdy7xa14m7va/8GtXdwaKWakq0ic3Fzkglt5FlxrvLKSEB8+NBN3h4Cqaz5cNwBL1ehzZtge
R4RbR+wZu22uYnMxdhOryALKiJ6t2SiskDvS21Y04zaAFSm2+mHtqZmqFk8wzGXeZOvf08FeszZM
aybNGUhk2+yBbzLsLd2YTIemkeuW9KCDWj9I1V8P9Swo+d7QZRM38Uzt6kNzqSx8OPxIop2+HvH5
sICQo9223kRGjrF45lml8yTpNP9x/F3hITINnClR2Mml6I6ekp37QhMnDX+Ff9zh8QUEH+WB7kSB
VqiOUXbZCGVJ9arrTQakM9OlIt3IO3SBehd2hkKmpdgKl2KRW5n2hk0gC0/KvEK/aidGieCxvaUO
md3VkZQ5ciBHAqa+3gnlXJ83U5Cy3Xp/jsfJ6UaLdgmSlLKgDKwFuMn2eFKBATA7siFfPpoSbtso
0gUiJ/XU0WygHElHtSJ/nvkjlR+tEJe1Nq+bVZ0+VHbeLwHGqukNTpMjlX2qLbeaEDLa1XoG3QWe
a1bbRRzJz5P9wQjXQjse4ypDGeLI9OWUeX3feLa5URvlC1SiQAYY5O0NaTB2CcBakrNi3UweTRnf
IxFdVJTCcLeivXMhxEellHE3RSMZSYwbmvcr3rDdTXtAd51xvnmoDd1CF2r8h+QHeb0/4OkAjnaA
qy+Ejc3E7D5zTP1zzxi511qzg39Ms895pzBiqahobtSqZn8Gb7qRi7Jtlqxod0Ow3KNgAkVmGbDk
zClshHBtZKl12lTnDPGTKqxpw6i7dewv56k9Xd7vazMg2shgDPnv08eHQ5Q0Ej1aGQ1WGkASYx84
9xE10xXR8fpZ4iPctmLbejrfm02CZdnFKKHCFFOyEL7I+DQrswv5U6ycVmXZvgNt4lOB/ruw6Fps
iKapOxFIigsgYYCxThwhHIxxI78N8fIe+QoaCsRBq1/lZvupR0A3LtjXeakgIhIvIkJMEYj0HV4B
SdFod92dEpF11TYSLVplsurD3W+Lh3T7mj96kI/RU6To8jFLjtMCwA1OO2r31SvRRVd8u62xu1r6
x2Z59klZBuKN0WkIhx+Nb7u9Ibs9D1rOFI/Rb+DAv2Vfc3FSJkH3cjIThdKS5VErPdl0WlAxwlH4
2pCEstq7KLy/ISWrd1/9xVktueeLzyCESlTsQBs/AfSs7AvTRq6wpf8v8C7TNgCZ7nOZjCbjMdNO
WR7PiGnUujjW2cVPPfwtUtojb23LgzX0naZna51k5qyj1Z3jMOH+uviylrFJYSwSDTYyHMJk0Vzc
cGEMyJ5CDmxciz2jmAW9tzuWC4V1y7sEkDAxPvMRs+eYKm1Ha20BgVtE2MM2hAq13QZwkLiH02rs
JcIJ2KD8S/PlYYCqXsy/H860mdVAUEgueOZlu4PWDvDUPyvlTvFiyuqI5HOdsT8cuUPW2Gcr41X9
KhfmUScZjIelyCaegkwZgMUzP7TdL0t75OrpQboF/JC59v21G9ee6ILwnSrvsx46t/lDeiHaHt6a
wm2lX5ELjXlFpPL6GMNMhjvSBve7YCN9fqm/kHH979yi/wODBno15eBbvh97zpyhOyUpT/d0MBdE
wM6JcTa05yNXA5DFF7OwbWhIIAsDXaSZqtus+aW9TBtJTPaV7Zhb1Iw9Lkpg4ZBohWRRQ2stVbeF
Prv19s7PizyI5yTcq/9Otd9ZiliqJXYpNyLzHAJQo7ZZmeu/ukpUQxuA6GUGN5A6Vsa+2EuiLJA8
tZjOfJvx/8+36+aGUe0bfSiYQzfp7fGiKM7fHrVec+cdLT8/O3i4V5oTtswmIN1dyPYheVSt8Y+Y
nCctoURbmvfuSUJfJNx5yxPGbW7VSwYb79BfalfbebFHKDlVCkc+6+GbsDbEp3M7z7nPAudHRJ3b
s94dkOItLZN1Q/Z1bHMPEFY9uhIJ3e3Sjl4wIpLEnHox8/u662ssc0rM3PfWygZFLic5FAO6o/pK
1IC3oeeYYeY1UoTLtHBu6cnvQYXkmanQUoUxEOXcyhIlRZ5/0SYVks2mgnwg6GoKKRnMR3WKOfFI
S0uAPbyMC66ieuZbpcbliqk9fQ9KnSF219fxSMz2xK0e/ED1WRp7OnIA3gERcyORjiKhYa+7u4GX
LTUxuZbtM/vI/t+dL8Q4zEfY4ltHZK98mNjhJ5g8YmqHBaBAd1TRwwA0ZjFweKJ+wdkIwR5Lz+s9
0jU3kllkQlQV56nnx7Qa6P2Gr4EGVtH3HZseGv2txxmdwA6sQoxUaQfBcUFHtvu/XA9vQSynrWl8
+vbppFhfW9DJqpzOhzvJYTCaH5gsbp+kmehvyxklcozb4+UR7gCmqZll8uY3jvS2LDmB5lscESHI
0MYD+/8GGETi2wdZobGMwnzGLxoLjpBwdvrGNRHuz9Eu0SKrogVNGR6jhIaCPbQqtjR7OHBOYEQO
0vHqngXDYZqGFgXDCARbBEQzsx7VkibYfIQ2YjlQg8iFwWKzbcHum20gaVozT83gpqTObMWx7o4b
aCwQZB7rcmyMuIbLT4kxziv3QgfnAEOGUYAUpcb2iKL2I5YALyrIm/vELPiKiStDfIV3i1FA62Ny
UrkS0TuoCuVUYjOjqPMNaNxaRyJocvJuF6kttWqhb5KjRLHTwqDrgI+wywr2gGZZRQWLKwe0Qdzs
B0n1PF3u6LW0df+FWOTinAOJhN/WdIjm/hCwLciIGm4bAZLy/dL0UYkjOnoNY3Ozn3eMKT6e/eKp
skQ4VV6SBWPkUwqBaI30DmJ3kR0TVqXP322yDN/vL3+nbnKn0KmXOtuOZI/Qwn9qRYb2A3ADPdMm
8I/TaSx7CdlVFRl2AuOKieutIErdQvCWl5cZ2FupotFc+BC7/A7/SplFdW4S0FEhrVSrgWzmlqFP
r5f1l6jkDId61HZT9ztEvj6mRtupYdLwoIpl3f8kEGkGNokzMFFy2xPmMIHsIkARnA1pbL+ZuIof
nwXLvzfaAk38qbS/cmfx8ueSlVt7urFbMAVDzonPS2T5Kq+Fpe4QYZ0QeDfOH5CK//gfmFx1Bs56
ixtvLxeKOTTOdzMYBW+lUGi7y0HA5MtwqjC9vB4SbnP5L0ZsWMvSsWwswx0XoDhKaad/YAp3S9F/
TE3zRkOUqYBgLTMg9UXKKYpOb4xQkqYItElAcQN6zHXsbe6Tbyu7McdRAr5jxP0mevCb/+Kjuwg8
1YREhpdl3hsmcqP+GskzA4fF2Ce30H5Siieahgv6W6Qg9B/AvK1Y8xXGGkvyxnQjWXr6oJa0nfK6
Lvv0l0Fvsr6HsS2WyVdb4Ue10nGDXFOva9zIjSysYtNkpkT0+/0ZkRiGIkP8M56mv3aF8mjFX9Lf
7TxDK9atPMXHU3VzvY7AV8UrQD36jOqNpopcUdl0TyiBtTdb2EkRYAiPxy1mNhCnBDSrQ1aHKq9w
8xHgjJecQK5dxyOe+4Fot4HN2TkqMKNkGmxyPrLB/wQzL8dkmBplZC2COZ7w81uLkW5bFdlLx8Mx
6PI0lJPizpglvm0KzkvKCM83WZBsaMQdssKOAnuWSZ9ssRpe5mNtEJeIwbzOOwrZovN7znh5ebi1
wxh3UfhO0/+jO00Vpcr7JCV3lk579vYn9bYHg8tLF+nYCKd4IGydwDcBBj8F3CRSvRM7U5+7rI3p
wwYXEjoMn0YbbqufnUvpJDt+M6BhzcwfQdVMTATzCx3jGAZTht1s+yxm/pZAskV+aoZKP4dn/meY
uLd9PBmqx9m+6JMJI7nHqhVLkjtl0WCA+PX0+82ksds4nFKoSAY/Nvb4zsjRe9Y9PTbeSTs4OGUH
pRx/Th+neVmuvubM6OgSiEo76Z3MjG0CtSmzwZTWRI+11fDbzkvUSNGGHCQYxowZ8o51CltJVVyU
ZM1RjIDgCEYDr8AV46CFfJSkP2/BeVRJpMXQZy3x6Rrrccok6jvT78Op9QYbSzWBGNbSKF2xuaDX
fJYWC+5MJIigN8P4ZxaL+l6/vBoV675KdLfjnfrefRZdpVZIRV8yFnaWVy8W+RfutZlmmsnppAbD
qYi886zZuvmGbV8i/GPS2w0pA0bF5bC5zveU6KcJFThWA+aW/JnyPqocwCrPz9WV3wXUDi8cHMlz
KbWVn1/SgmjyjIQMOy1uC29BB9Z9jh+5fT4CZVG4xazPKyOMX6BY9h4pSS0TFZa/GaxWp9JQRoX1
Z0pnzk8bXSwXC/qXXw0ZaxbeDB1AwQ+DQd4YbsCpJBuWeyj/jA6GCn9YkI394BJ1f+rESUq2BDWq
P17600s2QJf0ImJJmmWBdtuim2j/wS0Pv20HUBOlYpt0CxRfYsWc+8KP01CY/vUycEoQkXK2Eiwx
lp3sNGfNhAP0UIWKGQ9HEVzCIUMQKfpDw8qSSCTLpUKVSS/LVxLvm74cHQwXDyK1Ofa26z2H6AZM
1+M9GzLH6nlcpJ+4Bmu5SwqIzXXXkFr73kxH0pYBifv5qdHnRO1KxYu/nbYfDooO1ZoUYjfz1zFt
ojexgHEkoiMaPL9j5XzZD+b8J4SQf/PTNZ0TVhrsuNhwEN0ff9aCsV9pesvUk7Wr5J6jZqxxLBly
OQHdJKPZKRYJ0iqppRA551MLcvndEaz3rfweVBcBN6Raq3ivLDoGW2Y+IWmuQnYjtH/5o6Uv+T69
gwI4mUpC4lQiSYN6z2nriGTxwIyn5pXJ/ATTyjUNCFeGPZcE7gH2bhuzC0vfN3VxGPYF4cmW2LMu
+gc7x9YG5Ax0cIvTNKvxmP/+KEgOl/c7AqAnLD1o5m9c8p2r11+ZNZsop/60IhZeDPhIDYDe0Haw
2vj9nidU9wL2O9dHLndEKwkk4GBzXAHIfg861zWSDpIIO42MvVFrFXPXBdWRcBYk5a1EFI2jIXLf
111ycrgXiSRb9zno43Fpgg++G0qNSTtFgZ40qEKXG/Fd2Y0c13oy468Mn+k3ROMhB/WCpveh3gcs
NEDAMwCYmG1nzNcsFP1gQjmeBGK9kwet2iykGLkhGcHAHeqsXGr/7p2dd/cyZzpfcJnV991LUTF+
MFgr4nzYhMUnPuKcIE4ivWEPJrGvxzc5VnR41G0e+WGroJZ8exxfrBMjbHz5tQZ44ts9gikT/1nt
XOvPfTOQ3MltOQFXlGxdqVcq5ZsyBo3v5HizE5rhdtYPbA8ey1pTDEuSkGtaCfxGqI9amSf4JRi/
nq5EThOwUklNP0KNxIJUArbV8IVzrbn7xO+r7eZW5QYyRzWDBKn2Qek7hOShe+A8qlCdKrpgner8
5NZVzsYZQ7GFphNIRvhfn73Rjbs03pORSwee0WSnVdtshJTJ5QwuL4kqZzQxOCOFD3Va6VDGn/L3
Y+fYpXjeCBAbYgFemw4pus/B5H4fGape0RkeH820H8KqG37iS4xMtZkmPS6WNgz4bp9TB+/JSwgg
u8FPiVOh5h9NnCF/+k5VEDpGks6ho5CUemN7guO0Z+Ispuz8oHnNtAwDOUTgNwuCWIJOymbHYWCq
sgZiIVMIuF1WfgMzNg0HMCWwhCFOtRQchb1s4hwD2oMuLWDbApbQ7PyYuO/MAeeo1Zm3FWd0WCd4
v8SGwq1dw0SbodLcqpTZJRuuat9Qp5V7duJhHrHwhM+3q3zd/pKVDJxKAMggfFNsxaqRV98e1sxE
qJ9T9RuD4HoB2WBdAHh0T3KrBqSPkE5AU3Z9sopkuAxW2Igkcd+9RP5A++8ZXoLWjtsEoA7JZPnr
qJT+xgNWkkwN/NKU6zGvricefmmD6HlW7Qz0RsYCn7965lVhLgYZ0pRHhrVLbJ/plbPPbXqnkG8W
EgD8fQdBnSrTknUQaaqYB18KEKmE65hSurgS+NPLZ5nDDxlW469O/GkXTi8spjLkvaKcuRtaVS06
GKwZgd9lhXDXNL6+FlcQRiAcsGoQkjg48QBxTx8ch0E7yXs0TfMVTTtd6TU/tzklZio/ykAi/LE/
cILCNnqUT1unAGS9MOIWQe37EIPnqNGuTMHVkrW4PkICkxl6/tGkKWzPQ+QfIw4KiXNcsSmikAdc
T2kISpDqYwQRofszBPTuRJwprt6GzL/5aPNZpMpmK9bLe2nb72YB/mwpB4mJE1/1ElhJcCtHkj8d
8xkrADj/LAVVUPcGBDkXNvI2AxnJF/xuSAYOpiHa0Q+y5ORK0R7SZwhNnj5pex++s48acByrecpV
7OoaXL8A/ZLoweSRgXc7qowyzij02pVx8X4sC8YTBARO9mA7es1vI+jDlXKoIeHkkEkMGs/A+w6V
FSyKNwCBVNxf/mmLhiVv4DBAulPdaq0/sJ2I5djVKegtABBeWSsJ3y5ZIBHHjuJT4BoP+F+MgQJd
W1Bphisy6uC6YSG54AkmQhh6+2biN/zVkts+JX/wNYn7mkgHp6Ity6rnS8XLs6Uo1xA8UDyMxgeL
ip3f1T5WfIdZwdCufIC6WQrGjsE/DJ3gheJ1XaFdj+mVGoiydt5MdTYTve727Obd+cHEjZnE3Nd4
I5IgiOxFjeYpHt0MCr68HgmRQfVZVLJ6I1tJbnTKbau04AUrjHPAZsII0n58TmKTTGlCCVhms9Zz
1OAvuqxp+k7Tm7zsBJeZDHMal5CI8UoX1tpMpsh7HWLbkcPr3Tf/hh7ceEcetPy6+15x0IXoPxES
A/qYBn2CCX6MYg2LlMUtodgtWJpT0TslgwO/D6cw5uI+AsTdcJjimrkM/nL+pCDzTa41lw7Nxfct
ZFvfd6C+5q4ZV3d/3UjaEPmlMRacR4QT0lScF/yNARNhOO+plr3be7Z0Tg9UdUqzdGZTmDdiSkOU
mN5fWkq0TEtJwNOrueXKOVPIW33W8ZTRSRvE/m6SbBRIpllH/RC0wysWJesTi7+QNBPjmpNLMuII
3hugTfjv51wOp9AcQjVJdW1uVsXsNzPCDG8B/kbrEtK+6g42dxeGRQii1fTb6rIkSzwYFF1lulHI
l29GJ3JteOpDQJohrB7YMueNVMbqy1ZEo9fmgX+JbGP2VbmNam1GkP56lEsIzY1lFwVb9OJo5g2+
+bOqu8r08lNTZMWpVM1UcKzGMYAnCjLeFDn3P8HWa2wDju666o8FuTUEBu0OmCSljjUCLJMG30FT
MfoLGWJvg+BSB38/+ZwRGdwlr2KqEmROXjEt2/hP9WtbOSyqWEfuIIyJtNkTlr5XaAU7DR1xAEyn
El7JlekZzGPrM8beAVZYGrVZvlyY4zfKhe9isyK78kfGvuRUoc7gNdUbKDAx2FgdvdTSQMjgxQ5f
4APYWlFtgGAtfw8NV0JvTJVs7tO8LvVpfZcjweJHoiGZFm8XsmTMdCFYQp+PzcfguV4bj43y8cis
SRtBL9yBFHcQ2ehGSuqpIXecH042k3dCUPSLFkJ12/r9PuArjVYaD3bCagZ/V10dvn6cq6fHslL3
uWTVpCFh4zfLRAZh6HQy8ObIMLytRjaNZpgifskIypPCEKx8J75VV7oW4dziiiqUckC4Fasaxr8b
jbB8XJbrPpJxm8WwOvsq2XV/8x/j7UZmhwTfH/Rv9TvO7KoDljyqqEV+8UOrK0zBNerhqCnyDpGL
Yi4bnsZhRLlVu2ugkcz8TjpwKhXZukhgGuYOXiXdsVP8CL/2Vnx6DNixbWzBiyU+cdNgZSsvOX6t
QDXg6muHgAvzYIFAwj2QeOX8Y2C/XpGOx2Yl2Avs7j3ckaZl+YsAlhy6BTRnW+Dc4xWecctC9D+B
XFcdXMGtPIGTvd1owEF4I3SLfS4rr09lbbMsdj8uiyoqpHLu3KsITD3FvrHhZyAN2jXQbLwbVc1r
U2mwNdb/Hr3k52jw39JlEwgrYun85Kkb/SAU6JRuplwt7pW9x2pkb4t+FrAje4Ht6G4rm/w2fOf+
2LszDrOsglvPGhIOOhttjEfDUnO9maSCxqUw61tZZeC8i4GefI0MzDRO5ymAoNh7hQAcC6FRcD0X
esL3DwOolTLqz03y5vnPCsxITkKt9W0BeRkZ6R4be2S1B5ukiOXaRuVFztebDCCJQlW/g5SeQLNJ
linVRK3AhV+ISjtEMyy/udCoiLuBjHUYraFixOKQdjeReT7OIAzA/IIAHW+mm2Wt+nWw8pVOgYdy
uCXky2Gq3BKE5GD+IYyV8CdFmivIJYhFVOGgD3DI4DuyGa/CndiARg0qT7PuhVkaHFQt5tQGBPQt
oM3vN5MiDCKLm8E5okGlbo380K59ZN1AhAY6q4LMxls/Li6lntGnrxQL4T/Kj1BNHtBxE8Gqswli
um7FO+1KqakD3OaO8RjL7pycpQiX9dqNQScMsxtn0517Ph0Qwu+H5sSWoikN+v5HybPZsU0rEo6I
OYo1rPgHtGZ6Q7lUT4qtHvSSUkRGiEVXUIT4dLYo14ZCIPMX8zhEGaxGtiwm+1Fpw0A8jXm0IT3p
eMtujM0as9RzCPzYsgM0z5BJnl5mE3YTfcZBZCSv9lY5EFRH7j4Njp8j8FFbgK4ZWwdr0+DO2uIK
ke2j/7LXvcQ+utXitPf5NfDcwlTW0myr98SGEOzfzb4T6jl5CNv03o9nzxCwcbNGvyM/dYRvf6z5
DDtHIv5s0di5eZRdJIL5vjJ//mOBp3nsYwyg7jSudI7OQ69JNXHLNJaW8OX7mi2AlNuzl259zNWg
gxUEvpRliqVDs4lQem4HspOHSOca5ZB8am7Ntv0SmgA8gD7eHBhD65vlXSYY5UUbPpfmwFSUOcpX
GH/v485nf6JxfD8aSj+mvzMYHwuJQgaocqNe8PSP0JnB59EJWMJnoOZRN1QsJFSJ8aGaFq9qOlWI
beWEYhr9hgA4k/xOUpKHO1ZA7UBhJI5yiyYjJq9pXV50RRgRxsputwSiOEqg03g+wrIvKNUfJpWv
aflRe9sArZ0QFrdS6b/Ez6YKf6gjc24ndOliTDLz63j83ikkpnok+ea9psQ20Dp30UANrI/abUU0
B/lg1tMzNpvR8DTCJazuHahJA8JZe0DV3RRfwjpLqDegTNS12n6q9bctpi5gbJFJ81zUnQdRmUkz
9/FeEnQ35PNWBeCIsGfdX5drBJNlfBPGipicYUGRO8xBzHhyAFnFaV++74VAOHsxw+fFJyY0xvTj
46K3vAZNaAbQP+knqZFuYc4sdspKyjtMKdpdu/iRmqKtB6qUbW4AnMd9xU7arXzpiEF98SBWhctw
/A0Yxu/riprJ1S5PWZ/FqUae8cIpJ4JxfE/7ZrFSeKtVvgJxKnfhUHMnXrNYBwkLedaOcZl2DZeo
knKMAHFm7zBEJfCwWnKS8meNpzjbao8gGii5fSZZKaafXiRoxCDdAqQzipGvZ88dxq+LiU11az4C
HkEKQdC2IBYATAFNdOwppVwrQnupDcxBrbcH1jDMrFd8ndy4dT1rY7rPfCXLYdprt8wBGNlwBIMz
3CwLf9ngUtkVyTOOMdPvVU4iTHrZ0JWPmKzoKGDCaIO/jtr3Cy7X1MTr8tuPWPkWbLPejL0HnmdG
ZZU6M9RoBD9QmzNU3aG1WzKfyNECyo5ghAsI2c7DWZ/M4Iki2ECKFlElFuudH+dzgAQrEWegO/Hg
9ilB0aclI0QvppQcs3F0AfhGSqA33ES5EFDpnzKR2egd/JkWLZ72D99EXTzldhTZHy7Rom7Adzdr
1O43YNXDKr+kzNjioi7IISpV7qoMQ+TVywgXGu7DouSsoRSv77GIjjvE8UJwPfPjLgu2BMvYpFq4
cJc0dleJ52R2TeT2uvxVtHgPBn+GayNcitsZrAVRO/90ek5KxK4R+VucAGkazyyf1oF5Uid6cA+I
0h9Ss5q1BKyQp8i02stXIPQJ33M96eD5bK6N2RIBTlZ3CxkJY8JU0I91la60wAzT7y7jB/IXGHu7
JhNxw2dqoqGmIuNxB6H3uLN9hXXPl7XUoxqPoDm5bvvd+1sU8pUtXyp7/sr6603wSu3C1S0HnfUk
d32mUAL2/bKDt7cnFnh26PTDNYuC3TApxy8u4jESC/T8I1j4bBwSL0WAVQeHTqOhFwKCtZ/9YmUg
zfxa0zO0tGxHjXimZQ6s6ueJVC+D9J3I4vYZfwvCXUXnMvbL/W8AAcxSic3V3MHIv1dAT9JhwAEB
0LSQAsnyjAJjlw+/NzqE0JzN1G1BF+rz2Ga1kx2KYOeagu3xR1YP8yfkwVzsy3b1VRWz7Iw5IRLu
LAMGbjSSQ1mvlzgqK6DfXyg2ZF6zfYeq3mySq9qcoRW8+9rii0SXum+eZUxzA7NgT+0dL/3PHM7Z
NVQAQIriTlTZfj5UZmXox+jf0W9DkTyNZUrtOcL+/2ZCrQQOsxdO+bgDLUdx2/7SR2tvNhQkxSih
EfMAh9Ze75WKWLTmrRIfganfWboF17QrZxlPoqYEw/SyM1mrjaKyNU5vBWmCVoR2TurkzYsN4pyg
Kfz6d9Vv4dV9+00aLy+5JF5u+AmWtT42w7STq2cbZOA3MQ13cPeCb48S0iPLl64Tt3XouaEFq/8I
3vQc8i0btrfOtn+eOgBwmfw+ZtyNx+pmSM009YIRwmRmn/jt8zFZfW89Xrbz9Rsw6KqobrqO/vDi
maSAKlN0n7YZ2VojhCvPggx8ubmFrrupTOZO4aZ8wGLTRHgZ5cdq0gnEGNVBy7EuRx/AyRjxzmcd
1Ib58CLI81byoPGGAGbx3TwYv6b83edvOBmP3nze2EWuk4oP4yOUKicwPwUWs1ZrYhCDTOuaJBKE
cWNF3OCtGtOQSALkSm/hcnyCv6uQjF/FqO+gvyX7BiXbnWa737UWBdzKI4Oef5orM9MlDSlFTz5+
ZNe1zZXvTQmXAVa6HGUqQquRi/j04kauAhv1sObxX+EqnVD4tUPnG91nI+tjGYVEQzyoV8ZxykfG
ugbzUwM5/s+gbXSIioTuZN6aKLCJhwjfcLxUJ7o5a2kC23wMKlDALhTvt0jDLvjVipo6IBmO7Eow
YNcqAEciJ3F90ykvHwIyIg9bka2voR9T96t/rSVU5mBHKynVh733coYI2t3tjCPSGe+pX60McDz8
vr05L5n88dsl8wgxJUZXfLK2/WQEwbt6LEGjE5z8WNY5WapqT/Z9P6B5JJPsJpbmMoB4Hl1AQ10A
Pl/W1YVrHt9QMfExiD91MDRxcuAHs9PkmOSCv8xbfOcv4FFQzKQ/7CwuvPFesURKKGqC1Q9ppmuc
hC/lW9dAatqdwryH6DSlh6F8Z1uhvW1WYlczzYauv3gup1zKDiw8hEJeWyrNkrzZ/3uQHh5kwYmj
z3z1QhQz3R7+xxlkdrjJSZlUJiXlYuwAXeTdIO1YTpXZtPR/ndKq0S10Ow4BKqAs8hvR3o+MPINm
wv15bVgY4rpmSD/24Lfxb3rSF9ykrDCaiKYzxx9y75tM89/sqEWutP7Yfqp2MJsh+iT08tYDbDmt
bU+vxhg1ns0SoJMLjPx/v2HwRcA5GYZNdO9MDIe+CeQe7iXeYCA7ZHs3F2p6IUBObsvwr8BH/7cT
96VQxBHWhxQAjG3DmZ4eqaXI8mC1zDNg14gLJlbFfwr0eDqXOB+mPhKWHq4ri0FMOqvNAqq7Eqr6
G2+Hg7Id1E+K12l+9DUb36vWPevMRVaPDL7K7qQNyuRZMQM7H3YJI1IbPny4aKPti7E9UWFkfpdt
R+Y5J/v8Lb/XmD0rMGoCnjQx2m785kdFDws37yngCQrgh/Wp0IMbVeIiJjB8JD0QSJC9ck9+xizx
NUbwSxCtcuJzlG0FV1BIYW+9hONcJ7bNq1YHuFL04zu5UIVh2e4EllKNGRcxOLr3Z+iPVIsLtfr4
ckhzWQNK+iMg3KhblTQFjnOEnZFjvnPokNbLFbxVw1At4r4ZX1cBgef8F0JBbKzi2VxXX2fhy9Mu
DWqPn8a9EI9L2pbasQK8Q+vrYMZFi2lsdr9oWE/RtjD8KOvFQpYq/zurHwsU7uLEJaPkRL0PxI9A
Xdxum3L4zek8eCpPgoNfklHRTO4YqPiViuOWNVlra/OiPqsOO1lQ1GZ47OfmO1kN8msiD1IU+tn1
NWijMz8p7Fm3gPuUzZMmvT0d7gxg6nxiLl/6jvlDSl3qAhBiMnnUKe0U1r4TlD4yyFRVWxa02HAM
yGflzrWpA+i2jIhuZ3dCCWYyYmeQpon4uaKnaM7sY7/D6l61T2/lO7w/1lI2axTcuHJGW7L2phhj
gkQuOgvO830mn+O/qRtmb/riUDSX3w0zICKMz7YvVHOHzgVl6oBVNNoMswqqhRGlJftyre5V0o+a
QV3RirCcG2TXjtmi0yaWf8JuTSuO2bpBtEqiotU0O0C+feSRQGSwysvsarQ8lmMK3lXR/kqSe3XA
f/7oiKOOaF+mWuPPsY2+ubMZgqM7vS+AB18oibiVdG42I8eieRZTz9e4irdqstC4SMsZQP+NID7V
/vPVtIUmEly2UpFqHWakwfs4GJnZzKX12T2mItqi7SszHxV/8Gjt/KN67nzGi+3i0bzYyn2iHowD
WRPC5CzFQuKaA7skr28miDGzLpLUJNCZ2QxFJpIk3TJUDKC5Mi5cydl2rWJB5Hj2Oa38TADZ6oqI
IjH1aXuH+U7kradMw2xhSqaT+uJsUuh0896nt+H++MLpTgFiXYXUHtGyvJ1eZzaldkAhd9dT2tZr
Rdu7ziZ6iw6AevR5BeEFDFi2BmD2HT+C0wPbE/+hgZffZStDV67OxqbR/nsbpUcpMlX+AeOf4qvn
41HRHb8ABZkK86CO9iwfGQ3txS/0Gv1cbIjd6hRsWxJimKwQNKSfXbn0V/6oprTjmQrdEFSnBLyC
uO4gYrGaldd3MI4bFYN4YjdWtUU4dUgYQxLUSH17zy1LmpiHB0l7O55mjynHjDAkf/5BYzNLiZXe
8x5I7rUr0S3dhc8D+Qpr0L2CG/y6hudadXZZC9o83EKaoNynpzBDOfhDV9l/tqRmEEIgoih6fp2x
slvt8owflDkpRmQ3U2nDDSGO+p6jMZ6Z7J051fZY4rmA8pGe2WT+8zauUmQ8J/9cz5wn4skTiVjQ
L2gzVTT3Qicf3qc0YrouTkWDj9xF6/9gh+JZfXtfSuJd1PG52vMB31Cj6liAQ7UmZQreJyPIStBP
vj85LCr04hilCz4Ty7L67AmCNcC8GmYLgEm2Qt0xbYf8l0NYj0h2Lo2k1kVCPXLQ6xUccFUoJxde
U5R25CA/ruSxKtPev83ifnarrwRnm4RDHdicQ7t/0PhHI144HoA/SwCk5vBo1rcYFrYWQGq/Dqxv
MMZiMO999VBUYOl3vifzvSx8QeK4CBoURm5vOwIWS8/q82RLh3AK5SoU+d1gWfezUnGQbgMVRKt0
4tSkLVZQ4uhWy8JYb6AEGqvLaBwmuXVw8SJ5/YfVMAAIrfQsrgGiF6z47/A34v0Lss8VWyds1SBJ
KZnZADcz8xGzNM+I8BlKsQeKgOkdQ110REHfUZmDXVYDiyl2QLKFEuH0lHbGMjJwb2/FyMQNwigI
/bLEaopMbv8fkgGE47O7umA0+NW7G1eTXGFYUJQQU/eF2xAFNSINqzpSQi8fFflVFoj+AvaVlUVn
CE3ynoQJOytW7x1YhgAhjC+5yXX17xnxOJVA5DhmPlpKv5XflsGP8IropDAM4Ppo9KOaLBJ9eiXO
A/HF2FSGxVcs6OgGyNdLUVRSAa4SVfFCJDd4AKK2YUFe0jGoNVxt7OTTtxLbZ7jQdquWK5xjGBbX
+R3f7dvnF/a2IlXF1/9ArASqHdONeycOxAdBmci/4grox9oFJtMwUYHdy0ak1+HFq4VSgLh+mUuW
Waj7rDZcMa/xDlArKfhtsGVvnwHdCK5NxSvnSKjpQ7SICMohGMvyEnYVt0Dfe+ljmATHAF/W7MTl
pH9t2BB2A1AcNL+Ac065iJBnDkLPL14NLPIpt8VlJGBz5U+9ouxgUbn9FmOGpLte9V3ppKCfbg/7
ZrXNyVXPiiib6qQA/6DkHCiq5LchYxUZ9X2K17Ein7AFAl0FoB5zszCF8nBZM26nX54/yt0QtrHM
uPNXguMjt1tTYP3QqHm/HuyYnkSlVzdY9NTFitoxufPL6ZmGS3aNiXYxsskvyxsBXM9e7fCaTgfG
yP0JKAtj5blUcI7ppsYIm6R/WkilAlmiMde2tUJJM4rxjAGuShT9/elqf1++NOf+9vr48gRWjyQ2
kydAKzPq0BWdqg7cuvAWcL5+7iODlD9q/Kwb1/ulwgc2TtU0A6/AGlRap56/4pAkag4pqmN0+iZ/
4pQ18utkMSAzTa+ahmVMk7Hk4CWwKQ8/rOKSejB/5ejchzSvOV4dmDrisHLzl8OSxgGuSUiFQOez
ldFqfWH5sDQEyjbq2KdSGbRQDztLWkymJJ6cd3t+lRg7r1Hag8H074xEECKJ6xnxqK4zTSRhCBL6
BJUBo2+FFbeXW9Oa9mkQCUCrDOsk3JA4Ul4H03dYiT577LYpOLDKnkl4IOU2uFX4eG9f5WgYR9XX
jiu7XgovM2V32Uz12q3qx0o09uHjcsN6FEwV/ap8irMDAgMx4DnFloJZ2jdZu8kJR6dyX4XZlTrP
DYEujplPxO8IWlJ6wDdA2CYxWRMIsBrVRH0+gCLB2b8Mx2pyVj3kY9NfjyLGlE/5ETuLyilLvgjE
YAQw5WaT4CanzyZ8QXFbiotq4kqU80o3g4yLnqj8zr73LBthNIn4SFx2acB5PQTqCVO1w4u8vYNA
KD76w4+X7RxYg4GQWZV8a8/s4i34c4T3qiXErkTQUfySvBrVRadToqvDEgHgCiaZeAHvOdxdbTEG
RsHvU/2Mn3n4DIlg1YsIL6d7M5dFnO6iRoJWYBcJznkKQvAmptWWmNLSgp++F5TU9ug0gV2zAz8F
plisyTfnW6MirVn0FzLHMiUGGB6oNUTTi1cGA7wZxS9dEat34vELd71DdGBHrgNJfddS8ifksADw
+polOAps28JlT2ARW7uhr2unlyTEhY4KUgWlmUFmTjHyxoGoYQLjnV8mlXhSSmIEs5qIDPsfAWx9
eY4iwQkgliEeyse2Hua9DvnnDnuoxoDXCnRGB12ke+raWV/AcGMFPGQAxN1tkZYQlwT2lpXM7BYt
l3jIXwvuduZ7EgZ1q0A32Lhq5uLb1GTApkKyeLSyBz40B8l8x4gD8dFz6hObpgScqPQqfBY0nfGI
0rH8nXuipq5usReNBndwd6gcKeQ0YtZkOjtrgeFNNMPDy770sCXGs/M3VROa6xpjMHtv0k1ZYmUS
6x2GFNtZb8iwRCZK3DBQBNaPYLh8mxMuimYA0K+oNYby1+zMfJ/8a6fxG/RvU310v9ahDwi6vvma
iLP2qMZIvgOVt3VPUh0lOF2zLkUM0T1W8bTtFNIXvv8+/tK0DtaVbfwflRPjBtsYNJC+ug+DM7Y+
tRnQAqYM3oR2prCAFhOx3AJul3Xpgar5LGLhwqYrdVOLKxPhgVztTCQi6XVvNSgUPMrLF3tGkTsG
e54v6HSWEJW/HlX07TDXvzldT8xeTgC3EyV9Ld4PL2+eaMq1+8sSF0ZvfZ4CLjvjJVl6clTZ2YA3
yq19C2le2dxTDV9jcZSa8KrjiuRpl9Yml/OYs7iR/GrLujZpp30TmTL3KPW4pg0yDdhV6lVoxg3a
FCOVcR/ozRKPqv6Q+oKxBOEPfMebi4NUQtuJduDqpu6bLU53LwB3rWHe0q16+9knY9Er66u5flbW
K8+efGO3c4cBwgGo2QQvnnjsGOUlxtWPo5MA01T/606sFWBLCm/LqNXRIm51fRbAc+zNHley9HLx
Pol5zl/VUrSJ9G90Zk9iLWsRHH6/hP7eyYR043LD3PBb9DST38/sPNxFtuW7tATd0sQxLJmF8y3Z
uDIn/o+5Cg9dg6RUqFcuR6V484O3lwydlzkY0JJhxWRYW44tAj5gpfSRHI/3c15t8cRL8rajuwl3
aEEYLX8IG7dh4Pl1HI5QXqZfSrg5bTKF4GFnQREnFeMDHxV38ExO1Qqg2uykAlIMy3z7zD5dv6hJ
/DbsZvaUybY4ZbSWEYdvAsugZkFlaONTwiZ8dySQzT3keI9EV6I5uz6vJr7GPbs+zB72OOVz34eC
bwiGKTdwDCnyVHtm+5HaLfFIwXRv4WeL4htA+Q3mMdbecRiA5E87RGIRNnJphieI3tCdoJ80eaHu
skAhI28WLagL/mEHkcCbITp6dtkU7yAq3j81OqmTKutlQAtFWOawt6m0GKAlP+X3f/SrHmuyffVr
Io1JAq/OJXr3IZmk4MsV0hB6pU4KRZfuTZWYP06BP/UV13IRpd8fGTzMtjqGVyhtjBPtbkkuQxy8
iV1wErHmOTPNSbzBaCVfli+Ie2DAoOOUvEqogixnJTxIEME1/Biymn1A1e0+Z9ZYyrdWMYtFuotF
hrbN7sOUJ8C3qk2cdeqTnsmVlibKEqBIt8anzBBiV/JqhLzGJu6pLSaYh8WIaIZuYq5ZtjEzNz1H
dtyP9VHSgRsQCxZVpisLbkegHBq7OHLQLBCZz7HkH45tmU/RQCOo7jqMT8fQARkqv0p79WkdGaTQ
UWQ1SatUtXLXHSltn3neXhISiG2um7Twx2KPZ3D8MyaQozV3ZD6/7pbphgoNEWgwo0UmuLt7hpjw
vEhHi5tUiCzPKJ5MCvzoe8+sAZQwAP8tT1cdR0MTcU4YI4opDEUoO1e7DfotXaLj6HwAbp8XIDI9
AZqoThJUgvyKXueCqnTLkbUZjv8WL02kLbzGNhsuiLgkWQ5t+KXsdGX1q34OnH1d9mGD4gLxuNzh
5ZFbMSrlWB/eERSEOaakRmO3tUgDcPaZlow+pxUhSmWBQ7KxfjIppzydaSZuot1wGqUR8fd3lYSL
AB42IQhvW0LiUUHJdcHYwGjf0ZFi5lKyIhMTI++fROyZt2lOtM8SYf4lrMNHABG2/R2qTPsKUqqm
OKD+o1ont0ry0aNiPvfyE1xM0/shX7OnzQPHf8UKCr7jSdtLRmeNoX1fGiCx38VEjWzUvmjs5wqM
CNnUsokTsGcLH9k48/+iDwPqXzMelJINdHYeqBFkWfF56zecvevRBOzjqpTywUESQPuZCMeJ1+jP
IDFpU+5wPYld/yJaHHG8lzKPbH+kvyT96UTjh1AszSpKIcxOEIuSV4EDqnP6nepaBmh3U9PXbXlm
GDOIqCd6+X0RAFxIF38a1OLzWNuj37gWvrhnmfu6+hHSdUo7gRVEKq0rBryg6kuQfp6vedrkJmzZ
4W8Stt8QKHzEOwcmxEOAoCaCVbP966Zahq05LQJv2+TODV2EXZ24PLSGjKQgVTp0n16PUD8jgqgK
ykk1cGeC2y5V8fGFS84Wo4h/62e552ieUSmb4uAwKh3oPfyy/bCJmlfJWfWWqugHyD1jbmys4o6b
wUQffxWyKjfiDce2DtIX4e3+2D4o3h/zfOqF/EKM2sOMiru08qr7aJWwaQwsH08H5SfQMTK6Hd5s
6zMbegKx8I5oFq6iROqDiBiw/jExOu86S0Kygf28G8MawBFXaeVVxHH+vV/UtjpQBf32dwIMBspm
9UPsE8ii1yWjlTSzA5hJa0fZHcqEW2eaiBHCIvmF31xMHU6zz8ig/7fDEOUxbMuFABMCaV4Ft63v
EMOZmfjcDD+zU/J+hNYt/1k4WF0BRhRnUNx+n5CPj28q+jqLkypXkivC4uiMsBas5DJ/ynv+luJ7
Ot+KD3Lgva6w8TVl8b8TD3xHimc2y9YKaBfLs+BEvOix50T5C35Ze2Inxn7ZtL9wTJhDDhLIkMhI
TBsJhH7opYtTLo9Fa+mfWwKhzK8/oEdIw2T0h2cCiQCQ9IDDkV4eVPNXqMcmpK7BHZvIfxsb67HX
ILqdJe1UeGWO6AW2M0B+rxvsCqnqwuEmyvjN8F7Cpgwig6J1mymGItvRJJGTKGQ3p3ul3+VQG3+V
xWx+ZnzFZ3TTXIG1i0BJgO1AwvwncWHlDHMOCdKZ1XUXxT5qs4gBvJtGUnYtTJve6DeRoNC+aGDw
VTnRznwyQGa9qnMq3GeBOPJFQhBOCqLZy4/LDxnlMMm4k8CdhQWnLCPLJe73cigl4LrPnmP86rqT
Z1/ZxS5Q8azWt5nnPqj4Cqn21LyZKbIDl+qzcT2rtWMWt8/cu6/ORYomInQbZ3UgErLfv50GI+ah
pm9HX+OKZYFybDQXswGVMSPf3ZkMjwU7WEERMDMtucxVu92DyivYEIlXzFfwVtgd+9lAqIs/6YDP
mD6rWqdwksv32cbnbBtPjSsk+0llKtnhy4lXLSX0ZdDC4hpBhpgUsdOFRxy7vakNfWS27KULqAdH
+LjkuEtSJpD+knSe4DL4qVNoc6vQ7ICxu0k+cla8acSzdtZi+sdJ6rXknL1O+enzIM6HFPAHGhYm
kKRfmGxUO3Li1dDW6kUouauTWZd/4QLBqHxY3YL46o0DkWvUwVT8rjDOC4VMURhtF+ly+jiVGx4F
hxrojNI2lVesa3aybjKtz0x+g16Z8s4FX3IcMMyTDFAV6wbfTiNSF+YTQ/WImJ0dNlahd+PjLRiP
vna9bKYjFE2SfVr0gZZ/eqfR7JMUv9wCHEHlwbm7RlSK/0dQpXp3nkvquoRG8WSUMEA3GRUPjC73
LUdknUSZd6w6J1KYzlWdKeKWpmKra+V8VM+KJ1HxGky+pWkpoS/P/ehlZIbhV69utHUWOaa2l6gu
2wNv+2T9NZEw7ltKsKjz+Cto0HTS58cBr7Ib+Vqh9fR0fd5XuxhgrHL7cKiUgJIxjMGuDhHxNVSw
QHkyRntQ5ezazKVzKM69prMhS9A05QlUpfQe5pYI+T6FYfQCqGk2TJqJlu3kYHP4Ku/kswxUT6/4
HB9LdwQ0vacy8uITkdVC49SOkr4nJjPNZN74ljoLO7YWx4xMgWOcYLGNgWPvOE2qe/L1rtAF7Dfd
5gGV1Xb0e9m9dxkAiXUqfnFC57khsbLNZxv0xnYW+JdNMkkSUpDqudiQckcHFxToG5Rvm+TlFlS6
p8NxyMMDY+oskuJI6IPeJSmV0MgNc+Er3Ys7aaTAB+nN3t06t8lahmvJ66gUxBRHpQg6iYxNGXbG
TmZmSYqVugUT7hmvCQ7vbtAevomzmtGf4F0FVjjEOVAmdu2UiDdbEyy4mFT8w6drJixvh3RmGox/
vM30eeX8/UGmE8x2JpkjqNAxuOmoI8Tf8966x1fBDm7/gtem/enYiC7urc5tBhnLy816wpivv2hE
vHs+N+uhZ0DRvBNy0epGyg3uqlBZk6x9o+qQcWyjBQlDWNVwKU4uEwA4DDTjngoS197LaJiHwR+O
lTfP0CHxKHX73ncVjqUU7c58RF5vXjwsR6VpSUYSZAt5UeBKn4kl1NwzNcCXXK+wNWoxeir+PxV2
/dBN1Y38pvbcuUhhIegVjTfPgkusHSNNGEAJsixIEIRSqL6ruOX1Kd9yqQjYTT9Pg0nc14CEOBgg
UJmROppI9SIP3/Y1kK708NGXsQSTyVSs74z6hEf/j+uwyyTOLmWxaxUOkSoKcMB0mHmU4ZdF6Ote
6sUiXZYI7rbP+jXPZDb81tN1uze3tvfY38g3qX2bcF/fRfZqFBEeuusvbluItpTIEa4806E1z3En
zg4kVmQm8xDLq+G/4K3jz6ugxGPUGlSkemJMIdDqT7PmViHqOww/ywY+0jLZP9CvAplUVwcpCBHM
3Bex5OKH/AsHg4Z8m6e/2BK95axXYj6XE+WKMf+9FYhjpPwl61gbeF4tOeFNEVdMtop64MkOiIbm
spKillfgxIRrp7T7VOuPYnXP2u2Y4EiFUdEBqGdCI+vnezzx+pF7xhz62c06bhWTiC+I2IX9mCUR
pc8Vm35dEab40feiVWpOLburWjb8+8P2rAC3VkTM6bziOC0pXIVErvapZUTxtNdpbQsHNffJGiuP
OU/iVoTHhYvCXea40tAomv7xHGMWuM/Cx8wtVk/U2lCeM08j7KNq+6OreGFQYFYls1tDLU5lKzbY
/aRZWSBBGct2nLgxsWPuE+Ok17xWFG0gAGnKws48yaBhKgZbSKGN46GZSN4dxxLeOkU+6ELBiEWx
M+3P6A0X7lOfg5kEI2AT+Sw/peDPhq2Zz1uxB6+H+J9N1GsFjQUmjrIwEUfNbNpFWL/sEDn4dU/j
ZBSTIOGBzGzUjKXj/q7WlcCCOxYHpSBDpXdtxcNGM74KU8d4FI4vmu6CasD3KT0EHNAVgq7EzieT
JAcH8MEF+uc3Fg4wRYX4gYua4bjB4/hUsB1b+d8N/+KbDeudj2dfUQN6on+rnR8OTGsNdMe4bCa5
B6bvEUmYXKGTJf023VKwUYurjNP0y8zQtqe47bKMg+4QbftWSUBzzj3YnUCG+YCsDnkhqoGFi3xV
MXIPcJU+SSehHvSmmpOBoR99ZVe7Rr4NdR+6GROFNLqFuUD9MlhXAfG4iKnLLQWniHI8J09czVYz
A+HorfdfEn9uSf1Dcqo9einjgEqtKQ7fArC1q5lTsOskUoneSOyqoWeGGLphDVKEJob9XgkSFjCH
qBcxGy1tvyvmIDEH/lZzI+3UBv8xcpJdCaSTk5n4zG3mBF77LA/nBQ4tsrl5rLK2kh894WKv7oCk
QxyUMBnu/WLjDHFZuNTPiJUYXgX793+e1UsxSD7XThSp+k1I166GNTmXF8a7zpxFlZqukagCtAo0
eTRHHAxJWvcHTCBYQyqZe0U0dWn+iXap8Xg0bfYoZjMra3JbQr7npLuEQCVCrmjVxuXW0C908ccs
UT5K7LVL39wuRxquG/9BBG0e1Sdt/XhdFCU+K0/44jW1tEdoOo5+XsOnkiXvwpl1rA/k9eVBNZUH
8Yf+s9a2IVXHNaMDnKhJTrDP2TK3Qo2JwLaqlSLuZ+y4fnPFtlQst9TpOi/BrejCIOymUZMGQYJA
zEl07JD/Yf3D1/9sUnPeq1SV23D5dpqBCCX/MkYGPmQjrAA6xMJ1eAgcXiEj14xYXRUnY0PkVXD8
7F27zZk1EEjZDfZGfri/4WVY9GGah2BE12CDCi82iZ3p4eD2wk4LAzaSmrq0olPqKEOgXIRCvjN/
7nTvxkA+2I1pXg3V48oVFkf0r8iaypTrrung2grxHZUXyQ/m96xMi+SVIbNxhOzgt1L+zPpMvlrU
kzzccwO9ZaRftIoksjLmst1QGG/EmPRT9mosrNRdQiCofG5aPhqPCCExUqpDKoKuCStGi0IoFmju
scIF1hh6DXSwc/dEqqI/bgl4lgq1tBVMHvWwWmtdrZxe1C5qHSQkcjtLgyDp/D0VfGAOGu6w6ARs
hNHL1pSiz18j29sSDqwV/XHfPbRaWq/4sjEiyIfFPQ14fbthJvnMPrXHaWGUrGAe5kKzRtw9Mu1y
8uneNgDRVKgt8Mh2cAc5J3plInBdwj6BYrY1s+wqWNAuyMVFUQNJcagip9NABqgeYyfmWzuFOS/K
G1W106sYTBQ6gWbEZGGEPMkp5q8NAUQuu8dl812Pe8y+5oQFTR15o0dtrhmpbV0p/ij6h3tOuyzB
stH+KO2G4ivYbrSDV8nzljKqdnr4VbRrIux6n2KNc8RWULuw6Cqw+0RbCIHn4Cw7G0PfJpsCXSp8
wcDtggvA9oMZkkWFvSxim8HZly14W1c9k+yfASr9/NMelZDwkbP78QyZE89TgstRO31Q+5J9o3DP
jYzYE3HB2AfKLyZMpHMPPssPXCxs/MPHsTJRylRwO7RrkM+zaPUhSbZ3UiTimCqwQeUrWP4bycdj
OP0FiH5pUQvnk7VC46n1GzOAQY6pypHHTPQHmh0TloVkPxVq8muvpb6/WzdugIJVmcUHJX1mLbxR
1LTx8iXBCACMpDeeOHEgdH8uQrhj53t1bzySlIizGOPmps6EJgtitjDCOV/zmaXnkWL9aPp9po/7
w6TO0HzjgolxhTJkM/HdYOj4kUkWttlcr/kO/O0taqss0b9mY7p1+KTXrWAGqKeSwgwTEME8CQ+j
lr6IwJZBf178KhnugjgilPVU/rwcdTPDJk/BBCaR3PP8xr0+broEls3umAKOb85ikBfvxeIZVc0L
KYc6uc7hg/coAhvesqmcmEy5NQUIEpN5qiL5enppmZVCD6i0bXcOQAytDYbbMgtoQcbT3/l4ZFdp
HDYhrfPjjIVZ84C8JW6f20N/6h1E1vIFNKYaJY2wNzzcstcJ0ps8UmEmcTyJIVXjoS+oIjckA0U+
Cxp+pThxjBe4jRMc+OZY8u0p0AFdKbDNrVNn4JvFc25awG7EmNjJgB+1UPr/09gpLjGD+RmFWoM1
kEE4Wgn+ZV6gvGCXnlyG7JkAdo0kjghSWz3xG7Q9lyn/ECiu5bKJDpvTMqcmLZCFkW1lxlhQMXSX
7cGajaB6aDFwOwmm3Gr+sqefwueHjujjfw/RJFEuobeiXoBJVFuhptSb7OzoI1AZcbvsCm7jAF39
ljx0m0x6u1jMuE6uY1ddpqOH+EkK0gmwy+OGpGaC7rbQd/4I8xvpY3QeB+ftiManQIOsgbdHs+yM
J5+BiFIM/Kv0YaW7urOfo+vBTbhc/VCCzS6+KbV8fI6F+dTOZuPnVrvWdKz28347pukE2MogMx9w
Xon5YkgkB+loUDdXCt2FdKBGQ/LDez3hVKiCm4iKWEC/TCBgmvjoaECSnH5MYW2UOPDELxruxN+6
05CpP7vc8rlap8GD13dlTe3Jx1haoocvKiVe1SDFm4MOn4+lG0KhSxUey3HESmKCxausNPHEh8qm
ku12j3d2ezr4cKLjsdGQZICy/3ZbpH6cY/kthj7rL9t4+GLKYV/4U2ktX+zAk7HAcpKA9DLUCXWm
wvXcpNOqRUbc4/V0hrZlXckSff8cULh0GSI466jZza2ubJpmwBNMQUFXWtOzKZx9mjMDI+llV/Ku
E7HvLFJtLgVw7GMWIbtarm9x4YwkOKdsJzOTT8LuxOY/Ixy6TFwDm3bDgb6Om6qg3YVEry5nEcOO
l7Sj8Js99C9PZll+HR/JkB1z3g7tecAf3yeOjN+v8ny9IC70NHNeXFyTWRb433TVSNbtvd547t7M
DIKpZH+U4ra4Xy/RKZb5QCy5myE+IZvmWxv0oZHtbrkbdr6uM6APheqLKmHDKy2WDMyRe5mCWcfV
aXY0FZUV2fw8smR3F5TnR3WuIqrYS2J3gmhrcRFK3+B1z/00BQSPgtp9zNa42FsM6OKJJdJabjKp
l/jPcu3iqZorup+VyvFtZ3PBSTV/xy6lFJLR6f1Krsa5Wwj4WhoUaXBsHjmRU0PKRuI9kGMiEq2I
0d/rQt+yt2RhdC006vZlwU/VdP0lIzhwFhuaSwG6DCjWsV1NRsSqY+OrWZdVhQlZj9vE0hzriznf
TLen2BynA6jzOv4Y7FHOyadTm/Q52TXbm15jekV7EM6n1rhFLrZ87JTOaRYeT2fMVeumnRZtBmsS
vJUjORANYfi1WvsI8wlG5F0HtDFa4Ia+gTCE/spi1QSx/Sw9tL/GGrHoKDBXd2kiRzn+zX1jTc+Z
BoHhg1R5/O/6h1z7TiEKXOj+E1tpo1CsfPEsa3Z1v3oz2Ily7lk9ogoC2E0HEyTL98zJVDDOV0Oq
rVNMT8wPRIIYkgoX5G9ieoGk8Ou7jETeoRCtF+FccGD5lYDXJSmG3ozQOuwpg2Y2R/Q0IgczKH/0
vOP5CYL62anKZf1seA0+0k7oLFPKUxBMcNxljZz03nNwFkbQWqoflOH/RK1fEWlXJQestmTC7s2q
vc4S8KDCe4TEtctaCVSsZDmhfsuJC4sZfTSQ7mUl/ehg1Ard3F5zgf19DHKXN8WtQWqIwtv+7AGw
cj0wutkEalK2OoGjTbwF1SXUT/IcRqJgy7vrBnN/SnOtuIgj2KDuUY57sSpqbaIzUO9+P6vdZEtN
aVv5PK+JTDJGSKChxT7v5FZZU2oYWibtom80NgOEx3RdOOodc1mSgH8thkyGnmygDFCwaHzvbvkD
8JLDm4h0FtVZ+QZmpmxUwdb/u1S+a7OpMtFyex/ZU/xIpyL8A9lLx9t/g1UH8STtvC6GjImQLpNx
vS3B4w74U7wHIx0pavTC2jYR4kBNUfJhOL9Y0WVUcJNNsWKeUZslTphzuprkRNgaeKUeZi0WXhz0
XKz6MwiZyGua308f0XdRU+XyunqiEMxN5onPO09jeK36+ApnsIQn3sW9uow0y4FhIF6dvphlmJ3d
BLDXFrzAFTFFaFn/mApIZT9xe5vlOnqfcog312YuPbYIrCU/k+vZ5G+sKMxVxn7FWBc4tVF9s5Ll
+SERDyFwO1GlyApHtYRjdid41kdW+0cZWkAjbALUIV/hRCSVwaLfHz9pVvPzZtlKNMZEy1/rbgSA
HWSneCRyQNlFPJ/0I6AEoU760uxr51BG1UbYk/mhWWioY178THWDxXvo3fK2QHUbCIWThDDNVgyW
DOODE70HnSNfNDXa9v3mLBJ8je/SvJo3z3RTigBCJb4fC4U6H53ioFW60NKxxMI8JrUyPwN5mKBi
D8NRUI0wlcOgjIrL5ActYenT09j5d7dZUcUfjg57e9uFgsel5UbgHqCPJYU3/4wbPaA0fFUNTLOF
sjU4+3s3TYGOpE/v4CE+Hjcs7vt5dDot5GtAwfU3w/TOJ4e6Hx4JbdmQfyL7VkFM34qySNHhY7kC
JIcPDh0OpfPJVEWTE3wMNhdUMb9UIy+3HSFqvFCsDlx5WgxFou4zZuVV1Sn/n+z1T+Ao7rOYvWbY
7Kaqtz5DAVnMSPvsq1qwpmtOjOAJGlkW1QWm7bdBBQSJs/RCnENIdJyxi3ARjw3DI9wNLCqwZfYo
e0P4FfMbCAZmA7Maw6pL+GDGl5LBlniPXd0tBK9lTY/MGW/bUkJOkmsFy27akYdWcms16o5sS3Po
yrS2CQKO7fExpYHQ6dFRX869fq0pPyTQwh62WZVNIsLgBiUS9c3UZMbmR9Ms2WQxvi/m9mM574UG
nH4ZmypICySLIDM6e40aD+tnfPyb8oaCoEy2AFVbvLTlUXsvZAJNg19N3k2J5twHWLrGZHlDn0/J
ceYj9Jo8PzJuxFYYiw+g5PbYCueo8CttpTfzm4C4xmjp0EGIGHqF5Da/r2niZc20EQwO7bWp8unY
R0k55ctxKZvjpv6W9PV1AdBYhQjk+Bq2ZJbp/LQMkSfCw367vq9lklYmF7hWd4Tw4RzjHZKsWL6+
s6s1KRRTZ32Tw9vbf5azDzFmgr45arKbmyGYmukM8ed35yCac/o3RgHMqug/xPXW54wtM/vb6jhu
XpyqenQQ95tt1OMh+G3z6Xta2/YU/xJPkgJ1nwu6LhUlX3jv1V2LroS86N3/6ntMuIZs2ZB0CIlG
ZAlSZtvR1q2jiNHjCmCU/aBYTU1UNEa9MepMROoK2K+spPaL/w2YJ73zy8DW+V5XBsO0qbutg5cM
zt8k7EnMCsMpUbr8BDMgg3qlWmkNg94gZC8h+mgPA2iuEQFHDfidGaDgHSS5U00rCnnu17TLFS4y
TLl0HF5X4d11XqvdLxJdp8YBx+7rK8nZgwqIoSWPBK3fQxPUKCBoO2R0dqd9yFUWCJQq3luMUoxn
TusUyWeQj/YVBVCn7Sr9tamWbw/Hiq6qTQWiTHybrhM54tDid6d5WtuqKRG1/WJopmRl+4KTvFUU
YAwIZYeg3KtR3tBtu84ncrFc1+mLqyYLehvgNyeaPmSK7vl4q2S2rGJwcnvsJEWlkPepggA/hnm0
FLt+3HZdYimDfgKoNzwLkT72AUG1W9k/vlXyT7rMFVoEyJwa5bf7CJSlgXi9PbBs79o/r51Nsdm+
szOEeAlKfvUE/uCoITpm/YQMFkEbnHS0tt7N8J74O8ZlOkLKoOjDvGVxt6qukrwlFl5xRXrDkghS
ODHIT3XOW8nPcDimiz3/PNzjZLfYXOhM7wodLAqxTPFbRCZ3ABScfXclU2BOKHb6UjRG3+CCTN4d
UCp5ih/lcOpjz6H8VGFBkhkrODNcdWhz1YjjWGdwacaj4AVPqed6It1Ep0+DmCbnH9E0RKPABCsm
O8r7FlOudVmjO9MgPDpMyYpg4yug2kqu+TJz1HNX508zIvv5Kg0ezjGBpokIEhwoq4yTGpl9p1OH
H13IqKUaSUpheZnkuRD9aHfg2x5+zf7kw6Gk+1x67LdfP7rbr4Tn28r3Yrt6uaTYK7eCamsTxUT2
q5YmbN94se5mhjmE4y56i1w1I6b4lcnEfp4lBc7USHhtZ9TUb4u/YXLHlg2fWHuopdSZFhA7hujA
i49GRshkY5VxEgkIE+B0FBdeToh9f4Uovu1fYVS7WGHoqW04ZbufykEmfEgx3YzWpCnfqQ5dxNL3
rvV+nVt6VHFK0dG9NUS5WldQLsYrp3nSVstNtXOR83wgyyXH+KDHthEb9nj3B8XqogQJ6A03ZTeO
oNRGyCTA4DsdUtQRsogl3M0snXqj9HQL9IajQk+gACLNdyROr5ts5A7UUP4wEvABqADSv1sn0YDB
RyvCgrc5fJ3kJ/q8yvTAG8YH0K1ZdMaU4mcei+DnDRhXAfRZTjwMV9+mURZiI9OlMyv4orwP9Ed1
/y0lal5zYbkFX8HUuhGIoHxHBRhLHb+V3SURFqCfsGsTT+ogbwjbaxXBK7O+ULCMLSWuFhWqcOVQ
CAAO9xfPSkJpK5CQxxLkAnIsQUoQPNusOpTI0PHrt7CJCuLt4heuhkmeO01ndzXYM21szQoHdzw9
hO9/rgf/F8rDVYvelI76gAiArcLb4WIrVyE977Z1k9czXVuzeZPMxzHqcOeoba9Sl/pIaIuDUiFr
3wa9V0AtW1lmk52Mksys8D+4xRJaKQuWmdNRqXr2bIxvhtZfKXks6lCT6aOjikIHlrlVO/2SJsvM
Kb/i+btKMmNJsDY3Hpf2SGtLFaRAJaQNrUJCzXXRPwkgfw5QYe6YO0Lv+FaDGJIeKahWCbppKoNA
tNEOzwJAbf7lt+OBPEwh97RmBf1X+Bl4xrrSP5EaDLGc+V5p8Z9f6Of8VOuQ0V7xnq8ZpkJ+dHnn
q2+gwHGE24WHH5UiI8VNu6xc2S9HY6LwHqdz1kKhq937w0t1XQQtuwBEQS+f2Wnjo3psqgIPnOAj
x9zmMpGggVbNBv0+XLcCUP++2JbWx3FdeTwbdlaiay0/cC4ZG1OCvDv06uALW774dBtqTE48iMCh
pvsDQkV/RgVI327g27w5ztACvcpyPsTqAgPe5ngNKpzj3fbJLS2AxJcAObRS+wduE/XpAtkaMUd6
2oyGqaCcCqRM9KhfnYbYmY88KN3qDJMTTO0+qhBqmEHPUkDnorwL+jdOuNC+piIloMvdYNsz5owt
2xXUei67DJfpDK2D5RVHFpIcEc1bduEG9fpdhcDstJiP7+zs1aYF9KIWe/RJ/Riq2qiN01vOiZii
I50fxB+UvFE6NkjUyFF5MCyWX+E9MOJSF8Nafc0Bdi29agC1ksn1tkuxFecdX/2UQPQ+3AcDj0Sd
9Ibl/mIyOxaf80L6Xp5pV51evQRiw/bUNcO+lWmiZuz98Y0djxPZP+zzKYZYGcxTu6cxN579MxXR
D8gWp7JyUU+QgxaEEjJjTCcBm2zqYx6vBXhpEOrzC3sfqbutB8i8bU3QznoDWWANg4tf5Pp5dQoa
+sFB404Ckh0qoX/tHyYVkL2qJmxIxvJvf3g6hYoRX2uexfvdc5s1QCqxGUQNwzyXh2GMBWeQxVZH
cd+VESPdRWqZ1doxoo0OXKfCSNli8fidRk/0krnIRXoGG+C/aTg15bFiI/ds0E3UZbz0sTLo7eeb
p6Phmz/TOs0Q6F+2FsH+KNOr5xL+/AmYaRVZwiR81J0N5aRjPYa81hZ0GbD2X9jtmLyuXdeTqtO1
04vSwaQqkwGWH/EhlEXoNd9F1uE1WjhKQJznVxw7+onB1h7aZ4h1M/+86OLGYnSUGZr5pm5t2sF1
vBM+cVxgpw5EWI3RIaFNx8ppqIp1iyLmIxs+Fy7OQZjBwL0KqKjkwFWOMmVpj6B4X7/N7z3hSkg2
RELKv/5Bpsp/r8v5ShoxGg6DyfRT6uvhntzp/MjW7k/LuBKYqcaZdfzdrW5Hf+2U7R5hCPGzOsHc
WUrXxqoXWc6AgItMxXyQ6kHlV6Z68WPLp0kydmh78wlnSfbc4qqbIu8LaG3OP9zj9k+OzJQXxSxo
91wpxmhrEwyzl0mW5zOId3qMWDMM+8bFskAC3aKeO8bQTTfMfP8HuxHus2efjz2r0EQoUKHGcTdI
xfvUPWNMi4xBcrlvSmn1zHLSZA/etNloDjJDOSC/Z89LiCh0xM9+xId4HSlPeF3+W+ZkKi++rKEk
+OHJ16t/4OIdDgv+jGdZ1rwD6iu/43bswLljxTsRrgoaZiwkxvu8j91S5wSdfG7pAOEhoSUX/vjx
vUc+UCcgpJaoLc/zpA03d+8xZP3Egi26cSwBwLDcfrYzpPC11ukb7+mG7Hj50J4iucXpqm5kx+uM
z0D8MmOEDRweV4kFcK5/7Y5Jc5ZBWtgRvh3HjR2pwNjY3leZKF7ZS11asCepKSfQpWuUav7ISDq2
oxAalhES2yTzsJ6otZi1dNI42Kl4kfwozt+LoYlHMml/Mv65/dKzdyOhq2qJDrKQcrTac03f8uvo
/QyQ8SDkv17wA73pIS2i1xdLivgLtDZ0d33WsypYS7FQ0wvcKx7/IDeDzhwWVWq3jazyD3Lg9hHP
QqcAwuUcnWQeGjFeITCRG/CY/W4WEuddDdlWT7vtGQBY5BEBAI3nRKst3jSv0Ek5exFbTE7b0Co9
GBf8XnUPX1YLGGMhY5ok5Sn7MfhExq5DAj/bQhx5XMUprNzY0Wa22GyBNLD7FnDoeDIpfZwii9Wc
HFtxAOgK4XqmAfV/SEAGlp9yQ0gI3DOHQM8L7WzPtmWD0PjRNdDEgUotw3DemO232cg0AuxCZ/aE
BfpjxL0Sl7unuFmU3/fDwI9PQt0LtjDDndWrme2kMBW+LjvI1LRogXOlpiRflSdhNINO2B/2Ta8M
6hnRSf0jXtFYkTZl1hNwPTzHaUC9RPSycc9nJlj9ZYiFdKmCwAolIQCzLtyocs5gMHYyFM8bRapQ
sx0Dq/wxyhwKO4cz33uaJyBAxvAgrOk5RHpoUHzIoPCAPqAbao6/z+CtMiuYh3hGPxkp7MynagCy
9ikzxL3Y43x0KVX1TAYjiVAlxdaf1CKxwlonMUMZU6J6efEf1pRTIc1Fs88Vut+Oadd1Y06YaU3M
mFUwMzRDPm2x7nNEyYnE+CeUBjksZFdriiQJEs0zU8VJXD6ecgIBRurC/f0QAdSJn2UbK0yS03AI
YvWHOOsQ7v/Y3ath3Dg7sEFJy9xtdM/yhnxaryQpdZu7Lwpv0+SdAS1PfDz8yA3k03dckgtLrE9z
anPHwWr0JM+YSMIVC22PeezAeNZHRBKD7XEEIt/X6YnMMDEVmFNdlARZD8uqC3XC8AzfVfrthfSz
JqWz4pfZC2ETcUzDOHMCbAcryPYUV2ZpXvJBDv2TdiME3qyszfW0VuTf1h2K9ks6cVeANa6R0A/V
RoQGDDcTOVI0QSCQHW7m9HjMVAa+unjj7Mz65Tin8K8jaVqTlzM+li7esAQrb6SintdVtaKD+kRV
K8uhTKIqvoV0jO+m7WCoCXvdfRg11SDy3tk4aLCA5zGLg0Acv+kkSrNd0jiitiGDPVidw+G2Tc6i
eAJfkble9R6p5EljLoRNaj9SfMB/XubTfTNNLeaxhuKVJE6X3mgq/USvPK8hiaflnXIzR2iw83OB
4uWyiz8kkkkaxuYYBP77CYtYawvInaknQ5OataclrbLbi2pTrnHwWkOjjj55qX4E02a4B+c+pFk2
i5Wgfe4jWAUmWnHtr46JxCj2Fg4j0eVH1sOr2kuB1gEkYqMcTwlDJ6P+XzMErxIswhqZqMiabXZD
chNu5psQw9YrE4SRzp5vDsdOWt99MXlZMCh/Sahtfi/84tpJ179s/Cgp2tRuOyjnCjsnSTgzNHqf
nDPRP0MegWn+G28H6lRjAQLVOE4g5vJBPa6S3FbEV7rH7wgNBUOhVLXidVCAx79x73cnye/SLmsk
FKH8SM+M2+dgPib6o2LpfYrNY4iuMrMPLgwjoIYo49rRAQwKjvAGxi176V/p7t2KmeJUs/ulhvt7
oIRx2ZSQOkhCfuc0LeA3f1GvcLKzy596rPEF7cBeRA2J+DK6E2IQjdKEgSYr4UZ9OWonW6S1NcMe
r4moieJ+1YhOJS+C+qQN7ZsFigLjVjzOYjmurdjYfCtOOHlx3DI9RE6ZuDbezdiWUXpEd6v8GV9r
QYDLdBGV8Lxch6LW8kiGO8sxuk0Gmu426elGji2aEQUeYbkB5bW6j8eawFEALreiHqrd7+m2Cfl5
PffpLyGAgPzjMSf5DW59TTNDqwKyymq6NZZrZfE2ZVPHwDnirt0CWyT7cOeO9AfyGmkiFdTTLwXB
YedzUBHLKhPr4RN2M14TTV5OWqjSLamComUs9hE4jiESbJlcaoOc0Ae8800SBV3j9jQDxw4rc3dT
/Bioup3YnwQChPtWgbYr7DqTsTWmUs+6dRpFRgcTi9sD7OqGCUHhB/KcwXMYsFdrpfDB4M/iszRT
P7nvbc0xBzhnVHnIqsw1hYJLs5lh7ucle1o5Mmg4S+muQVGRgqu7nYKDUtvqo/mONcC4RN1Uz2vO
rILLO/Jh8G+3EymWZ8oVSOPKCdUXKQGbyiZvGQKHY2ImKL7bTSK0JmHVDzExs5iRy1hE/Xs/VsLW
1yOSz2gixaLydon5ikW/Md4O2LpKhhVJWQZBFnJf5+zm+YsPCooX+/LJSOV/USwWZUPzuxcAXCP6
jGhYcHA9A0xnkNGcuz/7S/GKG19AlcMc3DlKy4mf284KeBS6D6SMxdu+zSfwcVj4PVqYCIa80kEB
wio6NtSJwH5fcm3u4JNPysVsq2w+XdofmL1LW+H9vD5rhF5r786oycy9WcugloDoYnyCG508zCKN
TYBq3nrd6L9nKUeChS9YYIkTEV8daeOz6r4tpYqkuuJ1QVjXRL44ZKOEGo78pjvs6c4HWUmP3vWP
3GXs9QUF9QvQSrhwDHxjOrHm2WrTCCtBekiGnV8XUiH0n9dxGVuQEWq0X02PSksM5x6Z8C7pwxYi
7IoQg3AcWsUd1auz/gseVTC6r260iFGoKhLyBr+SNmt9RG3AvPjtZ/NVX/BjbOv4lejEyWWTDUYw
FPQqJLFeWXQQhzYpU2kepHnd/EujhEKj9E9z4A17t2Y+Gi2RU+mmNVi177weoMVd4J8Y5odeGFJ+
zd4jHca0OGBktGPQu9mdceZ5JgyukJGyJeYr66jXUnQDqoDspZrk17RngzqPKfb+lOVEe8cpESYB
9HPL10adLU7tU/EFo8nd6+ZNwLOHOA/z1r80sYdmhTNLaRLYMu8A4yfVM6/h+ATQ6hZvUw9u2tGm
tObDCS7CPYN1lf9Kp7OQ9UAFHJkMASmeNSDMc7QXph+I/UOoXo7ssj205X+duQMDXrRUmWSV0P/d
fU87f1nZXJpU+/RBx8xQ1BhgB3QXXTScbNYbwlpUUsHBAZdkFKGpAHevugJZmYj17jwPyvfGqho8
nbSfK3qQG2WJdtHcTpQzqAUKL/qRT/GlGbD0EdkIID8s6tm3Kq1gLftxlexKaEYgqE2aM5K3WzRB
UdoWsm1ynbgDH0xfXrlTZv5l7RSduWM1FdauBX8Zm8VCGBk5oZwAwM3emAYvjRub2dtWfkDG1MEg
1WnSWp04KMSH+BAF/AApJQjH2zNL5tmbgfeJiD7EOloZ3jWYDdkCV5KXJMsxqc17vjkaY6Mfu0X8
JebP8ryph24VQyGGloPgeqvT1TXAKjEj90jHfRm5QRugneqPbpW2u/5kNXXedYxUlO24PRSPBWEi
gmhsztY/EKrKf/xX2g1xxQsbc4DXUe+rp7bVBzjVda6NDfodQuyS7/4L70W9VPIRWbjYt7UahA6V
NleFl3FdOdlnexRKiYKPp5SjdrDq3YuTF+8mZ941QZBE4UG89fvVSszRGp2akdTjzI+ylHTeT0Hd
vUP8uEAgFAmkbDsKF4JU+EUBRZQZGp94rW4RICWBWJ9xj9s4RNMDq665ePRdAFp/R3x86sTDBGim
FLcMlHio1R55pj+ooT08T1SFGp/U2jLs0EDxlEkOAYtiLAPsz8bQ0Pwt6AQcIOPKuUmNF0LKsUIK
WUNzdZdYUP3ElboUuB/+Gc+eBJVT1rRgdvVTi8cZ7u2YPb0y0QBL2k8wweh4JEwkLpKJV8GQWHDp
xBpBsEnHqZkt00rDLWHN/quUqbNXIXfGqZyktGaQZwYIvCsFwZq1CkmIqQYhMFHv7XxwJjrvhj0B
LgxXjTwBKoqqrQMrC2Css8/YwDdr2bUqwnN9JdsH0U6IKHPkYbh5OQPCZmtdpUl31C+KDaJgEcWU
/zh2kKWpFPMiFDeK8G/P7dMi3YOpB/DV4cFA4IOOvwjRE7BJ0WdfRc5fWZwLCqiJPNM52vDv3nvc
QaNQytgBvN2NpFfdIAM+VBKH0qavJrxHaR82VFikm1QOOyMKAUVLxUMjEwaZPzL1Noq/uLmqnZ81
Otuwyc2uvmWVSXl8mUBPYb5YnVXf7CdbDcAHvnWc7lVIYC59ImfCtipwr/RDUblUNOQZCSae5JuG
tE3iQsSuekM3x1hEEaFZAyLbMJGGT4mjJc07K+IhfUtlRzVwJVe2J0Dw5qjScrTWULXPKS0tABtk
0J54coOVkR59cJXm3hmA7hPxsyRWygrHWS3w1VfLVTQV5mSQmheu4aAyR7NqvEEN4nY8NY/R5ijt
2E/O8wm0rbkONzwpydprGLzhVxuxg76MxcCRgj/6AD8FolWnWCJotuAw6BHJFcUIJblbkQE6zRzL
w/h4a36SZNFUF85W6IQISxsU/HacPnY4SlwQfyK4sPqBIMn+mg0K7Nkkl1J8pnM+RlasqTXgVb+P
EGpOTsCfqapkY4uzuNYDXfMSSmn96vHY8Cc1sZePVFkwzK4VuLAkeGMdj8F+7MPEc08UkSfwMgrP
qihhU+nLe0bk4MBXGQHIZYubgFsjJdBuOGUmZPAjhoQWHmKmcH1WMKA+L357C73ckZ4zOlRrsbnn
4VZiJQa0ifC0bfjGM+opil0UuC5BwTCb8WJkVeyoF7a6QTy6X2IiSHoOZYWXDi8DwqVueqa/Q7lK
OUvq3/U8KBfIp/p1cqbWLPnWuUnCzWmAztSosMYi2mzc8ZdMppG5uxaPd6ZKIzfnKmj14dkMG5TG
HyWpB+MRDcht/UXMyKnue7CKS56NlRprLdOFP0Rc9nRaEr8spnvU1egfdwjEmk9i4ThSfkTcn0e2
dTO9j7AbN8vACiuz3HdREzrqhl0L+53cDjvuIpM2TlTLqJypdULPplmeNJEgvZfv9h3ABAcETSOj
pzvIDTFjazJh9usoHVpe+TosTfNwRhyX2VLV9rucEDch0NuukuKZXBq7tIR+45kSjdSKkOYIf4/K
VOmKBJd4ThKfZOrYae6qz+QvkNM7dMRDC71EXEngRu2ZE11PdG9nYNuYJPbSlQbGXaLRJnY7ax4W
eifmtDwJy0hbizk4xtyW+XDRjaRfcKjxzxsGFfq0qCnhtrYA56k+BkD+LwK903dtCkT6e9oI6JT2
PRUUKKi/0AK1gEhCjUOiwvMF/hKPUco/cy17WpFgG9dWo90ckixto2rC6n/dczwm94hgEryrb+hR
t+I/QNNmfq6jy/FziyKMackiiMqAaO0mhGR5TTfiJi9t5hiXgrE0VLblyo64XBwhyRwJPZaMWUhZ
lGDMdVQsw+F9f4vfVSRMFoqBWVwuvrGulMVjjUVft0mIe2Gru3bn5CgE04IypHVjmr7kbz5xirm7
jqplWiEcwKkoDPqwMazwqdEigsl3odblw0A6OmrpS0yc65KZ1QeJIiCP/ktr7jQFBXQHn9CtrPU0
GjFzNDC+AnIwyLTEBcoxuz8zpzvjBTKLXkaSLy1P/I7zF74KWlNmFXzo6WusYtCxs2eW3j/w8mzK
jV3JLv9+GGqiRVwRH/itV5PPzfyertQ9gX2QouWMY97cdm4lBeVXZn/hF1xyFb03TwB2ZUECqcf7
RK8xCS10c7sm6spJWutpUi/U1b7FjIGGpQooZylldNTon/FT/cLasKyPNzgpD7ajDnlLkCTa33eP
0fBV0/aGHRCd6Z+II+0XFRLzqd9vhu8smXwQug+YOcNnH2rryPH1LEYs8FGvNH0mZ2+c1cS+c6jJ
kUPcmfTVof0jcUqoamb4kH1AG9alUhQAo6jf2Cpf0uqWvFerkOrDRQI4l/OnzaZpa4w0MlHWBrly
Z/E8XQSUdmtt2b7dcR8+QZQ6Al4nYXLTjTn3nzTbjLc+vpWpVBbP5YQpoGMH1Oqfoh7crhwcnQme
H/6d+JeNT0Fi81M8aNTWMESrZEbTZLYVqVXuyZYBUD3Q2L0cDcWW1O6RbMD1uS5HwekB7Urd4F76
fW/cCzm+VCjhsGNviKuAE7uhNz/0LEw4tQa/snxqYZoXSJ6Bs2jKrc879SWTjCPi9YGKGRp96uTE
s+lBM/WfjLYIr7lTdQMs4d54SNeJFQVGXFgO46Zq+njQrTiO1d/6EouTQCh/QaF6f+8+sSft5eON
tjbY0t+wFtN9DpQxhpmPQ0fpOhW/hzkkNSYMaBpMPPh9crmWkDlhUuod3sHA2NYzDgGT7ZG81Sr/
/fqd11yJE44HHYzhr8yK3KXvEvhCRmQBC61odk2vxTWlnFRYbPTYBMVJz1QBHKR/vJjfr/1TBNcF
GHnOJQLYLjUegUH8k+S8uN2dHiITlYSNZEEyVwPjnW2/gPfwdAlRI7REGxBnmUZRGluot1+GJQ/G
RNEZsPom+AzTaK122F7Oy2MfrgvJpuPd3FQo8SG/6J6JkgwhfzA6QSkgZQyAEsucwt7QH21nLjEY
wK/SyuD0K6zF59foQ6UiWDpLepG+qFTsdgYQJ8ggXv8TUjXSrpR8X4U+Ccty9y+asx3410u5rezu
+Irt+nOnC8J7uHlgoi5kbYOXHCA4keUw9AhDnUH3YSqJGPFrVdFCGkMy0LhJ0z0uG5P66gRuLsr/
pHsks5vf7iHlr1NrIzRBA/m8VdJddtPwL+/7DT9KVJiWkKRjkfm2gBGc4MmCUmpZpnkETbqtDqbI
I75Vyeg9l+aK96YXtJMkcsTrSzGGJe5JDQHLdQGOPMKaJlA9IdzwhgIx80kEB3DjzzSkxRwmWLTB
xBrgtFQU3hNsL1CaXduAcKIvlGAfOAbaOjclOGJ9qLh2pYkErOFMiCt7KHBQX+Rx5S4dUD3B6KAz
CzFFwr2sibDIs7dqQkBpkjQ2utD90twVvH+tjL7W2mGgblr5aOr7dK6Y6wufQljew/L55t/FI0Hf
AfQy/QpIc52bMkPk4mu8DfkY9Ci2ahas3yQrXeGg5z2Q48JG8L4y9CYQ3/C5KlFKUEH/LcDF+xrK
oBSphPQve0oUIsdBHRD2Pgu+5pqD/xnaQeQxTeddiUtVliX+7X03gbWCAsXUxMT4FkUk5h1hJsyD
z1wXsQL3abUGG0RrAVEfRRegOX/dkcKcffP/HYPx7BaYK0VoyQfXYf8A0EvJOY0pbPvx8mRJ60OX
lwqsXIwzcIuehrFS+NS4mClu8GrqK/zaRejj1bSJSVDA1lhl9cW2FWT/gHFeqPTeNMx3Me9KJPD6
ufKuDT3SxaYtxPsVO/aMNQBnynAaZ/v2Sqi/C1u2+SVmypQf0mg/YvaobUBmo35n9AfRluNB/hy+
N+G0IaUUp5QasAzwl1uD/a0Kn6MB/WjS1MlvszZoz4jILnftP5JeoXAy/X8zHeH7anuGCwp3diiF
GHjf29nN+W7vjNZX9VVGaefJ+U2LJJ+UjqSMUW4B3b3o8T7VV8lH2UPoEye0z6+VK4FuBc7ZoCRp
976MUYSzkGFeVlYkrZHt6RAbXJkn3TrgX1+6r2efH5QNniT5ys0/SAr/I/v+NEoGasnE13rAUv9L
N15FL5PtiQuqiW53f8qG0tDJuz/C7M6n6z8Zv0PcnnQNx+ZswX86yJBganeBnThilBxCT0fsXgJp
p4D34IuWGHZLTo38mn8Te+cn8F9Tl6SEUpkqrQbFqxhYRuqbjfcb/CHTOTo/mAx1MBcB4V4z0dFK
c8Jty3qrvTZJELGLqzNUer1zAjv9PxK5jbwUHFwVbbsmJ4eAcQM18PlU5TCBWQD43feKuaz1DVVj
LnH46/9p4wEZ25OqgnIHP9X3sszybZdAuMMaLdLpw4jxYpb6tvWIGDRjsa/7mMAja0R88fvXBY4f
WKCIr6003NEAkGaJFOfZOGDeKdfR7tHFEmxltM3Wbhy1HZ1J3h2uyeUq9/xtWc9t9QAL6z4ITpBq
stLvyP+m+CCd5kbU7mnVn1Jn8I1K2m8YbJBiq+aJvn4sjIc7plSdFErX0n316CcaOsj2dgO4FVh6
Cxh+b698dkFbYt94Q9HJIWb0DOnt+24pRz7Ba/GgCL/5yWwyahrMCpJe5xECbLHRr1YRuRn7upsA
x56z5ryLMhSDalbAKpP3jvp8wB8f2m7gLk1DOn6QhpmfVwbvssAESIitY8hlfn7I9hT75IfCcBkv
bF+a1CPhVVW/ENqeH0t5ZBE2kRwlxGLdArUzzsb/dO7d9qGfa9/7Jbrt/3cw727DETbI5O6pvpVW
67KDCgU7pNAE9lSvefL1Q46Qve+HLBOyJSeVGyWu1lOoLcYONvDfpqxpokCtbVP2MDKPR62nRmcA
P2GvMmF8Cw2LnnhtvdXWuzqAhnehBFzZwnX/uBxQwdMOdo0nmSukvXiIchQ2fx4aUzXiVXNh9rSa
Jue2zCbzGGZcQwRlgQXSZ73tXttoshIHsBtT6swO0iCZbLbVlhe8J/0PZoyHrQfUbmUKxfWek/rW
qpx2YPPnh4gQ1Sh+Wqac+PiNxq1Fk0Ng7DKf5Ehnekllx5j4pE2goDDaWwseo3OXYVsjpT++1cxp
fCEyy7JivJ79LK5hYibn4V3vFvdtbTQo/JPLDJHxDolEU+NGFpeOky8PYI5mYBLscQ359jg1pOS5
SM4TCryH1vQcqBoqQrckwH/PXIIlHCXuY81eC9UbHHeq75W2yiYiQJH1IZtAX4qZvuJYtVbyiT97
1J6dOV79mSAJNblcRHVpD8DFxKQ+hoXxSJYMVXNPmkVpZKw+m1IU7Y9jgGeudF0MuVFDomCIf5kW
DUhPnQJ136rl1R+80I5t+x6BbCykIXtvqSkmX74mnMySG61PpoMSUnpU322ZIEQzCl4CGo9wRU2g
h6ocQEyOJUVlBpQL+05cBKMZ/UB7h6k9j5tYYk4bpd+LlTPAqsbt1byxm83aA3wYqz6e48dZZ1O7
egrqOhuhDG9eRAGkvgShKw4iosKHJbjJUN0fwQs1NX51141TSN8MQJbHNUUnkAh6AxgRPLMAew2g
e6xZkVSc2j/TKBz06owWpuABeU66bSE+QT8j/eVkyj6SE5iyW5Qfh96Mzthnm1RMyPmNGmFbQw8s
M6UrXHFmqHhUiH2uyovcGqUsgcVfpZiKv4OIkpLsDREmiRt53OaaJ0MJUyi4qa+R5+W94Y1HJ9jR
OGcER853DPiCNq0PmNdFarWp5zQRRbGPlgnuqwLiuKNfcgvFuTVaYQmUyrYE/zfshwjT+8dn23+V
SRCNQIDjt1gaj8wF1qpD6xmqOZkilvdwzyc4MDnWitae6yUNbDv4LNlPqNkszJTb8iT4EgGt51oT
0lLm9M91d0AsjpBKzloFTb0TKWUfk3Ya5wb7bT2mc00pMZCkjr8kJ8eU/Fwtlb9Qdmro31AXTdJu
pnUb+vsMkNBlu9n+l3wJPp7HuNI+OLTn7zpews8dlBNN9VuJq0hJ3d37R7QiA+NgyNg0D8W49UJ2
JTlPsMwbELlzaBaF1irExe+QoEPUCr4JvsNNOcNPrxc/ThW/tg/M750z1+rOrhsrdeNjYn6uanjC
veqmIOGUotkZyrpWmHqDvj6qqYs1il0h/nzEUSBIxbyFm+fsirqE906xaSAiSyDWfyHjYLHoYhj1
WOq9prUCCYUd2nCE6V0Eabk53Qrr3LyboZMjv1jP/6YX/dlB0bHbsR7VZm8aAmz+j9EbHTDy5kcy
HELQYv/43ZJ2/iNqH9T9+IbhlF2WZ9lEVJ4jQtjPPapv4ri7YFpR1mVLTduc7ekri3vxfNIjDoFz
M6OaMN3uqaublxvZILIJOIpNpxYCYYrrWL0SkoWTmb9DbVbDp9kEnM0jmwQFS/RhcL5Ow3QeJhGG
HECVHBTJVMy7D1A7ejvCCZNo7bgA6yMh/6XjEylpWE1fHO9ybOlW1TACpI1LGyGRydS6gJBT1kIK
pGqOlq5Ak+LRDOO6SRIwKimDnutBooW4FNcO2xiqG8BcWHXgcdEDqqF1B1CvgFPnNPM8EwqvGUPg
a06q9MpaHfFYl0xAf42DuLKG1GAUjwq1xTsQCtrz/jrm3ynAzwaEuD3xkouA0RQhfJgRFNSP8JVK
ugwopJw2ZGdSbU3E7r2QLpfY3lkUtUAJZm82BPRmHTMA3AIQoh2X1VgmBobV/OAEaRNfIzF8b0ua
pkdsNGVxdYI4PgauUxEM5La4JLK5F6B8+wb9DH6ZLyMdoEmDRt7wF2GEUb4cut2aASwJwjDsvSeX
mW9mM803cDImKiuB37ZuF2QCm0mpEr2ySIeNQbbHM4fnt5jPWJtfa/OvCQr0OlGmDbFrVxeNsu3l
7A2jvM2AmZozZ5UdklUyqJ1fYId3gq3pIoIfCjdyXV6KLcS6dcUhfxLHmr259EBfXSjIgYKZlMWi
41R87zUVu2876/mwKK8GgzydOx3XLIHuLHDIGjGIniGt+Op+Tqnk4mB2Jqx3ROr0gqFbehOdALFD
G7M4hZicyKUNSrIXpXTbS/J52/W3kSCqIR3WewweFlhCBLbDLOlnnW1XDIqoEK1uVzmTgjs4YvxW
41B2UVb5wl7BfbzDFEF79pAbwnHXsYRp2Yk/4KUjguWiCh3WTEA83nrz+jNYiveODkKM7VNhbTNM
EWzFvxEC6fvH43lZYsgo9cLlXg/fYSIZ/DVAtg+yQ43ro1Uu8uDIDE0Z4eAVyYO1APgrBaIU7gBI
sLlgePXjIR85f/Y8xA1oAHnyGVRZIn0paomK8G1mLFH8vZrWQgvpj9jwa8dGynhk1+0SvrHU4ki6
khf/T8n9d96oF0wnoE/sI8yceR+4CPmKhv8sPm8x3mZ1iiAtHRxc8P+rXlw2PCcg/+za0LK9BK3t
BzXddQEgFG7GH6o8JtytZISOYA544R9XBiu2TYo5ejJFO24q6quTmr8ra7nwVGoyrOskudkpISFn
LrWcXysvexGblYR4xDk3aCjogGTr3CJcgZfduWnreQaBWzmLusIUN8IYj2tJ0gK78zgmMX0HZxhV
RU8OuolS2QEqcwEomcAD5zfs7cbi/KtEgCh2yxkiz4CIVADmpy4i6AGwont4x43PUceA1vdjkToQ
PXTjtvk8QUjGX1EsWO2EXBimHZkesZYQ//cM487sETv6Hah5d51TCByx6Pl+4+LOzMjYvo9evbd4
2+dHlgO8yAGr9yuq1pQWXDnOaeIAQ/wBIkT3QPEaVjVYh5Mq/cpUjTzrWMboso4sQDwmOeQn5zny
LqLyJIeHylvFUrHqlP80jYmGYk2KzFzjOMgNOW8bxzLDLzBueEHD86sHppl/D0snN5IR8kp2k3Tk
CziR/PyGRKSztlm8N2eWgzumaZHwmRR36VGCcgujiJ3JtTclC1gzgtD5J606w1y3TahgAN6BKS94
2mBOTRCrwgux5LS/Y5B2v6NsgoG7D424S8bPCGsTcaffCVfjswCifzsNXLZfO4ZUCjxp+/9wVU63
tBnnO7gXmw7hSDyyvd1bI2/1+QshTRIMEMaWNI8O4mDCcjghSYg5dJ3dZxSxGPkrWUcLeALjAvv2
seyBs9s4dK6V42bhS4ccpvw7iQPZbTnG3HG05BbF+dx/jtqiL20xVjy/nGTYvbAups0BMzq1aUFN
1aKhG96/SKh7MKqcs8opkrs0gqKR6VpszMqGkT0qoRzfPhJowyCQgysXmNYo5OJ3m/2Cnito7oD0
i9RddOrRF5p3QHm18OFhauR4WyCPhQox2MGzykxLHanN4oEmlDqqRzB9fefW3q4zetbApyWRYH7m
nSgBkLEquf57twHYpxXeHZbrxtFbIznBOrMf3dxeNToZEQUU2CxbuYOwOOGx3OZNRM9kCrdU28BK
tr+KD6PIB11MdoC11J8SndBovZofPcq3YxeXulMqX+igl8oNY9OCxiVJS4s8OCWj/4NgNZp53rhs
a7jqFbo3eKq584Hxk82kVGcz2QeaCseCItIeHws6ZZzeLPxlX4hKl449Ipw9Luv9QaMlAM1DeU2e
wW4tCrBicdHZRyuNtYlBNH8De2JdX7MIxrw1FdYrJT4xjrM+W1BAmsY8jxtwDDCtb9D8U6P2ya3k
oFnFtk4WWlVzGDhIz6K9fOAZeXF68NR1mtcm7FOuJ4xgAUHcibF8BNNSvskCzgPUWQUrPWkFL8Sc
zGXURFER30huei9eiBoonMDCDnzDyYb+A5ydQ5UGrg0vxH89+tD6pbKGlhu5KbJ/5YoL5eHPwSPh
1PsSO1HBNkQRdePPHrxZSZPOfVgiuV6gfgOtCMyDPZ6gjAl4UncCT3BAgJIxPz5N2jS1tulm1Jf3
jcF0DuAIYrjlfHH3/24n2rJ+YtMdslWOimjBiKRIEJe/QstEivxNMM0zEehl9+/EgW3fVeH6YhsW
kxQgPgJrpGpP+INx/inbUiFlDDovQiK1zINKLdVKsZagcPuYoQoeQChSsfjmKWRLlEdP4cwqIKFw
pEF9JPgBSv4ePf+oRuV+omIpcIxqoWmxugKZ/F19wloTFD6NtniEZqFglz6ghhKDIbxcdrVQMnWM
gSicOYre9GTqDA5vjrLxPM4Z9EkF6GIS2LX559B86DVFWQzf7XLPCaKn2kG9tCStPXEhVspOOCMt
jNH/0UMkz13HM15jZQM/Q6beEc8b2APM9+ycxoYs1unBOHRp+FDBll22DMrZfRhKsq7KliJOq2nM
I5TQnNp2ZkWH00ZeiTlR2JKpAaKDRQ9q0ae9uKVuiz1yeHe0U6jBxwO1ajHBIIjJcYYlgatIbZyU
7mFXCwg4MkVXm23sPlDITmZA6Cj9Zlg7meClco6hVY6bMMZFJmPC2pO/BB1p8f3SoyHnC4vTK+Qz
S5nVqR5xxBfoYTemcYbNd1dM1ySVscZyb9U4S4VqowyFEEivHcEOo1pIhupTwa6RIaZqlpzOmjyW
jABPXefnd2f2AlQT1RGx6DGP9FVqhKU6uYAc0zT2GvoxUN/Hichdo4qfA5GFcledlRJVPZCWIlAY
ZjzkYFuq8QCVoEwufiyQeQb8urJeasofG686D1xfQellg2+5j3MQy23nPSXuju/skY2oYzYMW/7y
ynbyxwIO5l55CzkXP1dNuiYMjPY1dwC0yxfjWC2FEgHanDmW3gl4DJMnF9cMnG77wnAvuH4yUQvF
01YcsPafXmKpadWCSmUaqGRZF5aP6v3wx0obmy1128sUPbe9dnFfTskR+U1Gdg73HIGdb2zUcFT4
0LFYrcMnecYhuLI4Q3dcvh0EK4hi0MwdqeOfwY0/0vp5ULvYpBXc5Th+rv/EwHNY0/HhIjUfojEb
lHdUrViSD5jMJezphKVXa0pwSUk4wr9b/E59ktkzGGpvw9ZYn1EfZx36+aGS7T/F75V2mV9SYmvH
87ZmadAUulV63p7eHmViQnl0eezxuTN1yXSLrGDbyx6+xbzgeA8Mu3CDIhbRAPEqQJYbr2Vt7kuw
kfvILYHJq94qkdhWkE33Pk2IQXdG8YqngnF4GbNb2gvMn9Kh010EV7YrRVxav4fGP6GRkMte+yTO
uMLx8R+GsDj49Mx5Mcl+tlWUyfU/PoYqvN9wNkYQ/yIZEEkq5XzhamNM4K27ZBXcNdqNl1Iu5Wv2
VMiGEgfmNHsuCJqptNkbssuPU5IFYdF4DKYY9tjdonBoY+C88sjQd0M6+iKo4TrHY+wZZPL0I4RV
jG9HprrlzzlX9AuKwsNcklpz+OP7QCGCCNz1uuCvIDm3oPsADBmaERPQ2M+WLTAiOL1Lu2Iksu8p
1nFDroALF1XzZFWxVHaT8GEyruzcIhrTx8K/J4ytirAx7ZU5/khoNq4noebLzgWfaDIzwNhPcZR0
YYw955gBqmL0y+se+bsuXRC8Tb9JQQl5eHIuKijZr2B+p8vo4mH8cAW7KjLd2fggxMfZ4/D00tgn
mCvF1YvT9/g/q4qx/DrFLxbUcOAsYo99ywYYOVNhrXfPzT7K/RLmgUf+2R73CIxRwRtigD33QqpL
PH66kNiY/NKjBJx7yW+rc6ddr1PnRskUsN6+G0Lcfjo4pGyTrbPfYrQ/5wic7JIjZU1TxMJLM87R
+DZTmG/2GrDRN76EmRFLUfys2OPDnjQUTzcDygcmx7uvGn/qUSyu12tU3OW52VbxhEEEIkneNm5p
WJJo9L/TZMBddb5K6hqSn14vqCv2N9wAYrj8W+mcD51MeCFDX11gmFwCT3OIbLiPmqk/bQFBcemj
eULYl/0wvzoRTjMBLK4UhR/jZ5eQVbQ1YV99cGmj4aY4wDjg+3NIoRridtPBijFgTFLm9xokaRC1
NsXTNNISbMsEFveKgquDw6AEa/NMHhJnPiqwgAoejwpKU7DSozTqCLaL6ymH7h1iFg/MtXe4nWb2
fVwMt414JN8CWJoy3m11aFX3sOy9iGJMxUrdJC/GftwUeUt5oEJOBhGr6oY8KTabJB1WJS8gQ52T
MqiLraWREjReTblvfiWKmjpEY8LOmN0f23o01pctk3tfYmqwFsKi8xIGysWNAqW+txkx0QDvcQu4
heRx19q4iRVxMSfELZaiQ65a9zkb/1SC8UFq2TKkxED4wO7vNKMX+fKT8hnyzq6ds2CeyvBuy5PO
BQoxQjzaKitgLmsLVKEQELWAi9HYaEm+LKqd/NbGGRB+d5MoiFEIXYGxe/SW8eZMKnWwACn0JbBq
+48SzVfyBho0i+ORhBmHPFDYT1EVfA1FBmVa954bzJ6wlXbr87KLIYquyGZuMnfDUza9YwLC6fug
4P6DXVzwD7Qv2XkMCbBjJxPTnRZm/9gZUrGGsOQcch0XrExe7jWCh+ISvHGBE0ANEkNfkQ9rIsN1
e20HRl2dxuo+7hsh55b4CS6ih4UZsbbVyiwH/q5ugdb2saOkDZcnl3iPMsTueP/xFKknkGxXHnYk
XvciSqbBpLRPyzGUfoUvuFrfrKUoaKInmo+DqchqhQUM1oG3mPWP9mec+iBlhF1aQdIRfOy/j7XJ
RvBuilzLGIAOfSCmtJDEAYdX67uk+y/8/TThex8/rbEvVsvkdyLIc99afbtiDSEi1VwFsCeJenAH
RL+YZkdpioMPJejqVQqOfAuDhx1A5csNmQWULBjZj0PSt7QyQls0StCZhQ7Qy4n136qLTfBTQ1Tx
TWi1Wmj1tXw65fx0TLOGMO+Ch5gv+spRlHGiJ9rCA1hd2jtHAOmxWKs7bkY300CbAz0KKTdnpna6
nVk3bEXrFo/GZL8x8W96ExBp9yaMpVyhD0VERoWsTnDQvzg4HKt5E6jS6gSAcOHwXC8ZTk/ejgZB
JEfwMSvmwEHpR0Hd5UtiA9HMV8iLb9D8/4AxTsFl2pw2FHXeGrKcJ7pnVJmP+PVnRnz0Q4DHeJlY
prGcKRY5x9WSM6MbvMjPDK2BbnRP2tCW4bv7YanP+RhUb1rTtLs3RVRX65HphzyIJuPm2BotJPMF
27Nc2NjeXyPz8WTiTuMgtvM2VMU2pLs509FWRlFp0NnzUy57HIs27IUrl5q7awkBEDDjVNAZ3unI
8+SJ4iTbULPHefTVyDxAW6NseVE79oMBYh8AMTcsYLJKW7kdtC7tnXThIXAmUPDHHJnk5hTHnnFD
Or4lYVSIbXBaXmTkyizXoS8VnB2i+e56JqU47tkdWn+xTsedK/cgR98zQ+o5fvNEhhs1XEJ/9Gpz
g2V/WOkOUeHGvJmQRgRY9kIMwDKWpOBUFmgO3A29OSgyA00lmatOZTicsFweGq65TW/K5nd6o9uW
AfC1Orb/xNJ0LKytXuCezdFNU3UUE7mF0lP9vJHBPS2AUUd7GPDEFme6UjeMD7RPWhtf9JwYLDC0
8tmKVt5dso4QT8yzEtfLYTldmmjmFkatsTHlce7DCpPRlb3ZsPEjSa5AYiUYc42ABRI5JHkkn0I9
HDkp5zerfDBJplOTXcCS7fUWVjMgjX2kz4/E5J/3yZBK7F/cdMrM9X31auFjTG1qofSP+OcT+7fj
ytdoIyRRSg9Pk+QNnKkWCTdzFjJDyAnJbilepiMaFbYB84eJ/+t2fN91Og7ph0/yMPq0R6cHUNKo
RTqvwuBIPwx1bVWXWvMDyec8GGbf/zIEafg/qnknlzGx+v1FXoAwgBk1umMMz/asWmTaGSze+83C
FjxBwu7cO6svDlpNAqTuk2+1yCBbjUb2KqXulvj3ORKRhPeBE6Aa5hOCycSyL1ScnLVEukTg6bJC
gCVFqDSsQz4YhRd9lV7XltGU/IS1ANYUjwulXplEIwF7BzbbID40oyS9EUzeNuHs8hrbKcbBlewH
ZtA+hDTuEEUd47wEXhUD6i0tKxzCRw9qOoEjOAz4rOT8S39A358cC7n3nCLt4pdzghtv1u98tBm0
MtUqcw8R43Ejkz3ZeHz2rhY3s0Rs9f7DWqhMTCuO22keRTI7XyZYulNDMGuuuU5AawFpUDDkNJAn
oMMLjY1IKwu/mDaRwYdc+hYWkY6PWeZZFOTL+lFEvR+q3jUFfLq3D0u/MIQ4V/rafSNAeMtVt7w4
CQZmZldAm7aErejoMNjN8NlahsVEzmqafdnY/xrgQVhYyRYKLW8e0qTtL8/hIwRDjpMYt7yvjpof
i0xWtvQJOEtarMXOzvvfg/YfDUAiUEKV2G5Jg1uAKcakGUo0cPRlnMAWqX8NfPAep3z1HkTUIcL/
KDyGjuaSDzIn9koWx1mp2pGogemh01tEMWE49HVwJwybUlBSWGZC5Xda0mcHvdZWLRdik3hQPUex
JRlfvFkdfh9VX9b9P2DUctfWKxX3r3kmN+m0ZsbbN68fi9qzESP7pKljoChyha9IGmlXKz8d5709
XnDGPNfwhC17CJ7jwK4mItWp5+0ZLgZm8QO8tI5IK5UbgqKzVQr401J0EZE5rnDcbBL5QVLdegAK
33N86s4+VliTC5sgqRNiYmflUV0wFfEJQ3vy0Ai9LVvo4duM8oUrjY106xw7FDwsxKktVFEazyTP
P+Rr8jRjIzudCdRKD+GgTG+QTSwTeFQSUOUqrYmcexXDSIGFCvAyQUXXhK+rx3hKpm8fx4zBjGV+
j2BoLX4fUMOiMglrfYbBlkdvNOlsMPwSf3gmNcT5TJexC5gc99/RhoM7LVp8ES0lY5H/JilMvEPg
8REMIzy0XFBkDAv9NhtObPfpGxfqlDBiB8nYEchAtDMTT4AWgg7BqDyQOpxghLgFpG46QCmyLOto
jOKdMXR6udt2s4UE9xhPl0RLkgGIIUKtV7iXyDa7YLrwBBUIdfu30wRE1hxuFmwLKX/zBgUlo4aY
nwEb1T1oiumvoSa63eihC5K150ycKUqMpt2Sx5nvVnLwxzlP1xf/5fLK1DAsRpFcf4X0DRvMCoEY
iU1Fksj2+K1IMfbZw5bTiznSoel36G9KLjG01PDPBqgDGtRf5RaeNEHKqfhhujY32rPTecLgjEOb
CNlO/qhdKlfSHt5Teac9EjtZOZc1P6FhwrV5MZwFd+6+/7RG/LNYGQGVsBNK45GEfOzMwWaFFvCE
ZanDfWmb35IJwqXVGIqmn0Cqqgkp0cdXskGLyh/im3Mgu4+4shPlcqL8jlKRZbnrS6l96jVOMAIA
OMpV6bsN+CrlvfgEo1uOKXeNOKVAHLoJfzjAHYG1S+LIlNB2UNVG5kzfT5tQSDENa6KYcfdBoPwz
w6AsDnQA9RRLtiCedBwQ0psaEa6sP4FDtk/C7IOUwz4PZzPB1OunNWgLGkTYPBJiQedJDnwidKof
3uFtIkE/Q+MakjRvASuetpvHxn784/m/meVXiz6Iydet5fkIhCmAE+eHtKDgCi+cqTXlkxK/L/hd
Wd+aad5C3/w2OKlXkVvERqyPnwmENdALBJzMqGJb/D5p8zD/GL137XtSr0AWnjMSxWYZy5lC2MOE
bOU1axXqpVX8tdo/aGYljm9qzOi3YF3SBeaEYgHNJAqeHX2pRft6Cl0azYmi98AN/Mp32KtSoSD3
rHLArxTvwrBIdM4TSW2XSJtWkgVGO9eAyiNxdwC/KRoYZajh+Ai0UNEe0+10O5C5sKv5D/LZgUIL
FEW0VLrMTrNYHoK6n4qdmqjpHvwsMUkn+KmeCEWlkNuOKkVREdxWNjI+ADjaS/azhx3/o2O7g0Ix
riL06x+1EQi145H6rEJ6b2bS/Q6ecDiy9++u1t8nyN80EmcD9ENpzlE4Vj+rMSB3Zqn65WZT6/c9
vsEr8BkMICoYhZHn0smvNASRW3IEgHz2GDCTzmxltnzjJtvjVoCS/heQ1PgpvPlc0ANE5fiDOjUW
smoWSvwsu/FjtUX0GKgjeQnDFft4Z50hLlTZrAOQt9tW1lOp/OlSPckQGmWsgFOssRzwgY894v+X
EASvlqSNLRtjfxosguRo3VSa0vnrgeCudO8dSVewQa33GmdJTzbVRw+9XWWBWqCsHFGJxg2bnVUF
hjvUepmUcLQXVhOxT2603rN7l6EuKQV/qNGzTFM4bql8w5SQyJLEB817Bp7DPhYK6gkZqnC1WBWq
JndVLHqZKP7nR4ejfVRe4tomIZXNa6tpBCf9jef2Y9yoF1xjWFxirTntS+tbnix891OS9k7dAN6V
UUZRe/bZCd64ZLZe9b8kv42Mq2cqik/AVpenFqombEK/S+tn31wCy9VOWx1XRAKNgfAXl9nPIKaS
7zqsNk/o1HhGafufFzuyprjnArgboS3yRl0mX7eiuMUEC+MnO37+4Q306XTWFbjGfwut2SsroU8Y
3EvSIWTexi/4XadWkTt8zuZoSJDgKyXetdFKhM/YecoUHjxb/e84c5NIUryMIlR0CGLCZZfnBt/4
ZTraey/c0XVzByVgqfzY+Gu9Afy3TFF//6y29VSS1DmNCSK3Q+WxPSLg/ENLB8n69755iR/nrhmi
Sos9R/FcOjsKrqoLnQDpAiVGSpNr+Ke/Ilh9yQIe8k3Zf5fFqI2oxnYZ1vGkHFW2XqeOThGn+z3e
mTV3GJsDCywYlUmPYD9M81o5VVKHUs5oSumc1kXKSdrT0vqBFZfvk/YxcBF7mX2FmafEh2fSOUl3
GiWjC2B7c9e6TuOFgKrCmYTQz/sho6ni0KSvbe/Vnt5q5UGm3o1q9/WKYgzXuJf61mmeoK0avgGP
6cagmDBiBepjVk62AY+WcPdxBh+TK2dOmtMLC/nlMWdbJJq6X2mWTc8n7Vg0CWTKSRmfWpZyZlY1
ZrvNMHhEVRoSc0XB+PZ/33EA2isq6gpoz1J+BN/ysGd3vAxJajRqwUtMSLU4IbnXqCeqU09L7iJn
YdjQtcMZ+SrnRg4rP/3y2QaoBIB8kif9XT7C/pikCQ+hrsdg1Va+rK4z95PQTPMnaZ+NUE9ddc84
E4qDVQcrWXPe6QYBET5UI/r+L3CmvI8t67m9ZUdPaoGGyJBKRUWCgoTsw8TaGi13C+5Qv7zhrPHk
//H4JA4rqqo4zlhRSM/E1/04AVcr+YCbgJYd3pVvhI1XdKN8/nkgovdXrmCPfSyxsNoTn7oGKIZV
AvYO75choraxnMxaltuendvCsekxGv8rhqkVhhgkbLZoTEgDsgAICCXGEJT5lMGBaDbi51MqT0G+
vWPwwwzboIa8BcW4uMTPncKNbybx2Ep36jhHEKvvAS1IFK3lnSzPdZrGtiyeEahTSe1NeeD7tGpV
JZBktfS5GFFhQEX5ArJuf+qQM2GBUd0TX6P9gS2Yf6HmsFFX26P7piX3N+ugIZ+t6uYmwxHVtf2B
+jOWW6JFvDXFVkeNM9pv3t2mKNdDxpdeMF1mPsvZOZlMYUmgoG0ltOaPM4pYNcAUnDgeNLWYZrjm
Uh2ZvxuUIDj/UqZo/oOeHg56v5MaAnsSf2Q2XyNjnPQft+skrytpOZtV9CsXXJ10C/I93SCqRLU3
cZ/3/sr4S4a+t0A04WQGqPqEx2O79FCKIkhP3apTk0B5mq0T/WmSlx6WxC2CpfdvUSBqV5fCd46m
C0IixP3BBmQC3tfprcGxwwoeZEA25GjdMwxBlIaWgjjyZ/MCqXFdqE2E0unF6PD6qbSzFIKxFJ3c
gSRYCHgO8Tg6nNKhOthE8vuOR1MIRuT77URTiN9KInQjZgOCg/7AOv5TJj2mnQCl9pM/uMZC85S2
w1L6HwaVevgYmcTtIUvWY1757FLyWyMpwDvOIcFC2i8N6VOschN9fTfaDE+6bg5A5LdGDhsYPcyU
Rma0Bmq35kQNWipDBiUstExq3Tw6ZW5SzzofhiBmbsDfd6xWRe9ACn21MgLjFynP7sLoGUI1RypO
u+bP9u8kUUCJmwQwVdarAlI0tTW3jYQn8uphuQrLPBRWixC6KBWuTJUFSy+biJJAhNbvsHFGFiYz
81hYcHpae2tIqW/DbhyE06cXknVVW6bvskm54XNrhms78C7ceAbMuPJcC6Z6y2U9WE+GU58URmAv
kAg1JOIBFL0JmiN2/gWfHXz9dpel7eLZWZ7XPHqiQnkEN9I6xr4U9JyeIb+bJFPwHSTcBPEWm29k
OOZSt6+/LwPn07Va1Pj0rLhIxtw6D1atiSHRUnJVqKkPjMf5a4/M7hkcLXCZ1PaOyIjgHlJMjoFJ
pkrwcPku3sMx/s9afHVIxwoQzWCH6JE1B0BY4L07hmHlDF2cvlwi8QJWnZKkZGlmm9AsKzVCdLbo
q93rLPxYNf8x0M1nzdrqtlcjv/9LGjter9NZNDarW4dpUqqPdkIaO+WgelhBxHuB9RhMYwKuF7Fy
7BvduvZAwgyPX/jjjo9Q1Kx7zwyDgP4iH2fJKXAg20I7R9Nla5tH1uCu2a+AOxNVC+s94Cnqkoyy
7Nt1Mozvt6nAhMNlJATY4B2DkU7qh7ohiHTLsx96JPHMvT567K9jFrhHXRGXooeVbfL8FM3YUkht
0N6k8GmULUwv0WvwpDLX97+WZTVU7DSUSWjSTizcrQ02Q5vT1mPRJW02tRMebOVrDAC49sJXToZE
bNoO3NZRMX7f87fkAV+Bn98wU9yiJUFDopPdDpY56ibA3ILZ8aiJCNreoSM2CCoiUe4/LSkYRGn2
jffJnGpeQ+gvc3Jc/wczTirhOCO2OFiozvHKFtOBtwUonKTlVBlU2VP/hc42pKOPHQVafyw/R0y9
aAps4HI8bMYltciOWSiqEPAmQ1qFLAnlCaCHqUA3JuTHLiRvtZcl17DTIdVC/AQAW1vzkPrUAHcV
4Ba4YIvGA+sYvPwS/Z96PzKfC/oUXOWLayLPX0Ok0YubnPzOR3Y+evGBOunWKYtXRriM3HpOrHgP
+RmHUnOsKlmFBnz/o7ZTiXysqJ4Kb84XVzweWW3DfikXELlHeyYjCSYDw9jGMLwCzYNkGzjNCKbW
spDgIw2JKd+YxLCjx6D89XdgqrM7tGlEsqAdVwFHhqHMMUjgfauF+G92YeVZSloZvVegU/WHFnSQ
dZe5jdTX+aVXyNfEAgG9ZEgIOireI0rVfd2lANhvFyExvvGBE3+IhWCCR2O2gf+LNJsrpDOnTAyG
CsvCX4up9qBEp2pUo/nR2tQ+W+5C9AEI7Q8iB1GSrxnPKfK4fOm1NsXsKRGDqw2vNhb91KBjLkF2
mf3oOQ5V0BksZuE9f2zXV9W+Z2FGhkMzd8c9rOiMzulJexFuf6F+ZNLLbt7WTZRFhz1mA1s44Lqj
wN55ava90It4jFWV0YpZsS8WTHzB+mM0rB7w2tbc3DofUiViJ2Adm1jiCGEvl03Xb8wPkn6DOlTG
sDjtj3AH/4NN0OGepGIW017S+E0kBKkjHsoBVe3wYqMfDUPjQY0l2Am1ZyUwl9HHv/fXdatTddk4
TJix1j6aJLtlfwsKleyj2IzYvqm5TDUnGSYpHBXfPTnSjYM1JIqFDjFv1LHxmU61CXhDYdRTNwQY
oulspZNSxVaC7aU7n6LSvT0fGM3pw8EET0MGbIdA58IKrq/ihjZIkhYKDMUPHYkTR/rk1B0hkzgG
jlJhX5JH1pGMEl7k+GRk+OBcnxuFTKmVMyhn470A73Mv/ZyTsEYscp5xu60Yyawtp9exdnD2ST8R
7PpchlwEmpl7s7a5sT3uFGHuAYwUk4OMBC5HGpEPVCvpZCjlqrYYggpTV450n5z4dAH3ByyHHcte
bOD5ke9pA2VhAN/1Sb1agQ1uVtl7roVgwMoQRiFoh4cbubrgKEe0Ig2rzkxb2JR/MSa21L3Yxt/B
eo0WLvSDQ4x5Eb5VzE1tDuoAGbsmS2pUvO3rsvo1bYx278D/aCrfvzSW8mU90GUIF0qcwMZZp2N/
ELrc5xBbkwALh/rVKb2CA+eE/LgqzgMIPeQaDudGHypGXLbnqQBveUdyVZ8lW4t7JQgYBcsAvzY8
YgMi38mWSJjx8RvTn0vcR+mqhizz1t1eYUo15qa7i3NL8CFvZZ7lP77PZgjVhjZVlzk+nw70FJoe
Zvh6xn8LZ5uU6Gw4nuiG6DIlW/2+U0dMTDx+Vxp0a1hm3lAjtbI6ekL3FWtf/4tIJMm5elQDGfCN
vbaKS/4VkiUq7tIgzqhB37HDWDjtu/3q5ZWiA1ja9lb36Ht8CTaG2pL2v1l/K2aDWc3iSfx0a2Dc
2T2PTVAPJFcHOIjMxX5lA8qRNo58K3SrVVsItGLKKNvIMujnzMTLBF3nm4K03QCpLd+gH4ec3sda
RIfeZtoccg2dPLK06cTl1TTA4jxPxpqEEDzEcyJCjmQQw9cvZTkWQnn1gQiPFp9XGuTfOaKYZlqJ
FN/tppvT53gid5ZrGIlZV8UzbBU82um6xmG/hguuTILUXskezWxhHmiezPjBwqNC+YDqMQch6bE+
h1FFe+bAUkG4SsycW0mLljZC4qHy5otVX+d04DqcLBv9Ozb77+7WXBLWITB5x+nDkzWubhquoPEO
QGw0HqJZ8GEHFYi3Ubkk7gDNaHWeSbQxYeLaHbvO6+fIrqyPC/qdIl/vLUohOFfVZyH3KYg01iZh
dSTgJPtYLt4DRPT1MUZ4uGYWgKl1jyTHkwePC6ZGkmFYTkldjhDe9RVF+NgtsTM7jDWcFwZNIAfP
XA8HiGv0zZ7wZXecjmVyENq4Bb4XnM0mKVn4RsFs8oY5ShL7K69VQyEfgstQzSo4xjrzt5OwzT6m
V4t1YMq9h6YIPhRq0gFD10kmwcc1tdrTs1lmWbQcmk1fJfnVA4H/o2EKA/ud/+ijNgCP55dVtN5W
5zq1PayPrNzQTs0WbL7WqnUC82IMfIzigbRw2QI7w8d1nWdawfCc2XZPdJPVmfY+NSFiBznI4eFV
BozDsI8UA99HWVpOdFXNVQNWThBWCOHvK3+CVqpNstxBlVBYF9YckVAKky+q8KpCVobhxuJgN/vt
xiiPuPdEVt8QG137S0GX2duO4q6nXJX0bDGsl4psFC97f6itNqSlstSO+JT1QfIDlYIRiDPb07BS
6svzAs977THPEaO3wwMPaXv/XSh7+rrDZDbKtqjVkt9luqBChZOpXt2ntXZdTc1AC2y0JdcaDRfG
62xfy0r0VKoVmor6fbowbqjfuFz1iA2iT1ur3oQez0Jzb5FwJmhpLcmgWaP5h0Q5isrWo9M4Bdfh
og9Qx9BqJl83DmyJ5Bm40lTw4DNejP6x2JlXaZ/eDthi/OYBlPMLUMR9Y77+o1c4+wTTC26RTgmT
YzRNXsIcIk8alOb/aoxp47Zl0i4P1TdkLDtlB+XESeq+6FTAuG86zdioqBilkYT7uO9fsOBkd1TQ
2Df4TeSsJxUvHZYn+pZxJ6PCJr841nRboCWOr/zDZKjF+aFcWcYiJStBrkIT5qEp+xWa5I1EKhdy
nJE/IcZAePsY2tQLK3ZctRSKnV2pUddN7P43p6AxSDhFgihqW48lY6MHwnQjKegb0LF7DpIIacrg
65FnNj9sv03GHp6aBhV0PgSnNe+/0LGcrW1C4Wb6jelln9acNhhKIDkPLExG179QcW/io4hbwzWn
t3GZscMoACGHVTQSON9ykULWVluVukLatN4yLfgXnHXnmJgTWlz1Je/XZ2AVL4jcpWFMDIhb3pIS
jOZtr6z4kT0AoPkaFtbWKcatzRmShsovV4EAT/5EhlrKjvPzi9JgzSy4N0XHWh0JQ2F11qERuPiT
qhem00le9EdohD2r18D5aYKzDgeF2bpsTtW4/KmPxq5fDclx9en2u4vuPF3zuexwXHPfAoOqDqiE
8cbbsmk7n7jg9z5qLlesVJQdcoyG8HXleFWnec8NcIGdOWlgsMM7aUKildW9jzY8wdp7t92TULQD
CF/xVwc42dsucrYWZat4oyTr0//G14mprKHLToNwvVu8MN96AfNhbPWYcImc0nDKa35ofxEG5rh6
AXsjlwpaH+R6m7OK8Rt63pmFgSrxIXDXw76GPZ0OtgfEWaXH9vCpMQGNyi7Uu+EDYgPGtKlQQ2tY
V16SvRZugDEu7I0LWftqVscVlZVo/Y9fp6ph+ace487YSa3h8C+kOO6Ud+ErRNr1oKstNMNfMNdn
iQQa5cH27sDyP9pxPfmZLemZygq5/tJVofV0Aq8co2Vyq9GODMABUYvY2qzzzcJHSUz3yT/6x5d6
0Jp8ogqQFRO/iPF+Kr/Eai8wMk/bIqI3oVTW1hi9p+cu6rKUH7E7lygTY4/o7MHCax5XCyFWV28C
fJTx4iWVfe+gwLBOGV9cdW+BxEOldW8S8ffgQ28V7MaasZsXLCK9XytvPwStVDPPyqzG+vQ2VetZ
0FIfetRqY8NiD0HA4XqOshcHrdsfhye8EyhsVTMlFV5tVJLMHD0QF51Fkf1K1kdbqgl7MCOy6c9z
X1e9QBPYuivFAUW6VceoiEd7nR0/WBs59D+ODdiRy8NaxGQwgT6TIihYKLj6PhO6R62bHXHaj5+Z
MMrQE+z+zcYJYNchVtmwAoyCK8m0HSE8HKNBf4G+MkikPmd0awuRL5nXH0ZQPsbuJ3r5fLVu/rxv
Xbmf4cqgxVNtbuVEoTlpofsoOhePaoFhNQi1ZHaemYgvuvcb2UAUse12T3ggQsrN8gebFSKjbU/O
XSaACbyQo1IlQAzWY1+nXqgpJGK+VO7ecPiQRcMMTYioDPPpmei3IOHajV7+VcveCED6cGC62Z30
GmlpP8Z5/MhqDtwuJqhDwCb6cRC0DlB6LTFGpFG04TjGzdEaZSZRT/ZPQRExH//QBcneHEqzD2n7
ULrKCnlyqP+zqhI/AY9pKwHezWOQA9nowMoYYs8Bx8XoA/ufQMHrKHQ3i8rl9Ef0jHUdLF7KwK5S
yrL7sAaZaPovWdVqn/M1+u1qC7srSnhA7M7Pul83c40gF0y6jcbX4lhsjWEAtcxeq4DlvZ2PCovQ
4qlMwmgiE8iygsa0xC5XdorkF0fcb/CbUdSBurQGI+dm8fvoZWmYFKl5RiCeQ+uKFaJoDsa9B8ow
lwheE530tUFuQ25LkuDFC2sIPHj6s5gqK5Df7xfZEDhKWL/jaW10JTDTyrXN6O2crCo0rDgNtk7Q
d08iIr/MAyzmviQhsceU03cPlWMJfmsRsSUWtvqzB8eoTAtp93g0jOo8R2kkThjW57XRE11nBjSk
SpUB1qHVOJpOjysH4huuuwV/ZMiKAHSgS7pv38WILxRy9aewn+wDlN77Myk18Wbjo25K6e+l9FeU
cn51Z7nUuM+tuhu2OmQVd/VnaL3v+oECoo5fREByL0K3DaDssBBeDB2ChBo4+eRv5Ad1vCchax0e
PShEvcp0G1//snI0ImbLnB40gJLVks89yx1kZW1s382iDbvHIseDri1RH3jDy+qGCBHtcRWbPUHV
VsJKvaGHD+FUnODgNL5DITFFbHrC8CXiB/9yC5OPxnezT8kMOq/FLS6NpXBqibbqo5IbwiaX8UAa
8HFZp9z4/T2DHmb/BpTpPczHQhT0GmopJwp6rBS8Mc2oaw4vTlrqvfeFn6PpAorYQuZ5sW77hpdx
0X07OEK8qqDD35uDrbBEYSydl4CV392wWF7NmY1FudpJv0Do7rVaVG6CjaSDDTHOxj4S7WvvTz2d
kfCGQ60oJ1SobRYjkov13M2dufR6L6fc9as0JpGWyeAC9YdFaL9GoT7YwYDpuDkXthwYlymDPk4x
HDu4maDE+0f3xA6zc4AQSBaK3L4SmxvqWqDsNx9mX9sBG1oA9Rgp5llDPIIeeJu8JhzjLxOsw3j6
7YFx7xORhembWXq4UvG7YoNNw+dd/aGkAcURJOr12jturgubzMPV22GooY5D7KeD7bZquDI1HZ7E
uMDn0ykEasJv/D+VGPrHVvFrbha06xugVfA0R4INQ8MQoYhCu0uhWQIRjno2v6v8dC7auN3UVxVn
+JPAtXh8igZVw+2kwiE20kHP4CvBEhsEfrqK7mR7SjEJWnXWyKLgdSZ6cibLjFkbL4SSbcXNHskH
8kxSVbED/yTBZ8fe/Vrdwh8kL/uxtOhqQtqblNqseLf4nogHWCMlszePdRmW8hKNmRlNv02Dqxd+
PqJ1L1PgpNiFQUSUkX7c5o2LPihe51UuoNDE3iow8iCjH5b8kqit+TX06vf1ihE46aM3p30QLbnq
hGfh06nS/68QY65SuTg4DYfXEIhtDW5B+2YmgiOvZtb91QTZpy7wPIl/LDWYKVikFtWbSbqw+9Q0
grAv27vIYM7eEimC1BiGRO+YBqlIvgolAhQDR+o50ElWkAIjPpi7BWFee7IUQ5BfYMaR8pBsZHU7
xobUmMVwhG6f76mGIRcK0lnIkBH2XUMkZOCsBDpuuj6PLZx3Co2mdRXKrc1nK/Cc4wPznyoELBfT
fiqE3++9LGQe6aALiKZhrrT4/iqvucGHZ0RF3gcHK6Tm9qsgsV2hzZPOw39ugkxZXMSCRI2UFb+T
2e1XF/+P77mQCT58VJIRyrSsI1Q8/UfJxu1TaEpXe5+HOJ+daAESvMQZguDOK5yxWskvHDnkKUQa
k5Q4L28RH9ISdnWto9LpC/AoCwhSrsNtM60c1yMrbBdRME1zqs/MgKKFNBecSzEIjB4/5LjJEIxS
KRFv5ni8+PN5IuGbcR1MwTEqItP5seKnQYKdU2GWhnF4c7MdE1Vo+RivP/T407NKprBK6Oow3Gj8
gQXI6zl4/R9g1zXrJF+DKbzQncM91yPUE8vuYXQU5XZ0k4jcwvi2bjz7IViIMWEG2J50xuZHaOot
/Jy7HeKzBQ/7Q8N0P+/gwSTuMM1y7GuWDSuiaCpx8ZJ//kfYQzvVFK96PYbVMzwmqdgyqCBJ1LTN
dasikbS6Lqxs6W3kUwngt2OPK5SFNSyjEgMjMyKq+JBJQBiUfWP7MgkV/T0F+vgSOPxA7E/niLc/
XDTAoSBxBFbWrRu40kwXkzpArQlS9348k8KK8QJ/50/9n+7F7xjdpZwzVPe5oMz6PkhTC8wnF16c
/pzNBsx3doL7RwVAU8vhkTvv2Yyubmq/NUQHm0rie/PVgmbu+HEE5vYVoPi3DpBuz1Fl82U99caD
b4AJ4lX8qDlXX3i+P8zzLwFpbe2X0BuPVGyzluceQszYoAek2MXR8l2EqDveqtn7KDm24NMrsBwe
p7fbgjHvD/0xBhNlGeRp7a7r4TWpCvCuCBz7n7+qrWrXRjpyTuV36EzY1rTLboteQT61lJyDto4V
vpTS3E5KtlFaa7Mr+M+0tbKBWLnO1W8pagvTqcfuHKUfqMB2CrATdkC6pdKwdueRSwZZYFCMiCRc
AFXnCv9eXO2n1v31TlrqK+QmAcMuMiSVp0oQTzHlHhGVx21ZXWHIZKz5mHJAh5a/JfIPq3HCFbVq
irGel8hivIgSY4c2/KCPraJUO5Sggje1y99BLS71wm1LSfeXwz7KbekmJskz4FgU3zu1ld6yQGbP
F37Lpo5f+K1vTaoCnN6bgFh509Ad2Ek9gJ/Ij5ATVOup6zRQhkMI/NUAthCNLJOdgHtdCuzeZ7e3
P0axlsHghIthGbkYI3XNemHvT9meDgGafdeYhyOw10T0vQ8dX7MlXGts7YY041UDXMS1oUrDYUPK
ElNvRBMsAw/dBVRDSUv9fvXUj+aDbrPv6g05zP506dlQHdBq5PYZ7okQxzQcTG1E+TxIhNmqCytW
Z10kwk+86Jcb++OKIAdJZnBhA5LrQ2VGheqxSzuPLw18VPWSsapEA1UMjqy8Es4+d9n1d7KWkftG
t09fNczAUpBHaFd04TfSoRtfAqMTf18fFTVXKBtzmNp0ojk6foD4g6IKu25ba4IA53FRSM871OeH
jOMuyCc1ptkmGm/cwJ22ipbUenuMNkI5lTkZ8Rob/Unk6UJERzufd6BjTRa/knVftMarhc9hXxd+
KubyJXug/zz2aDGyKvTUpsMPzrV50Sv2MfCgY/3u3N8mV05aQ7yeYv153nFJPr10IuUDhCG9UFvR
fefTGARhB0HVNmIFVzDxYAXdW+CFEO+89UVEi3ilgtsIuEMCxAe2mdUiEOT/RpXMBmLIzwXr1feG
lwEKyITZBPm9Z2duff/mDMHWN7kZxv57jDFZwU+GqfdPOTprKzYm+7pgjRUqckKD1T6eZt01JRjt
faxK+57QPQ6YC6Sbv1bvzb1DPn6xXZBUoQ+LlCkldkzXgXwALfMXGQevkQ2c/4MSRxi9YVAmehT5
Ghjb1d3eTioucxx+Ry80p65X7oUtPpBQvg3jI9PrvmrT2d5FxQ9fXNlX+2zOOv/3yVvmyNodRxF6
OPChEMu1dAI5xfkAbMJC+buEH9LkhgPY0p609AQfVL3Zi5I6Ebp05Fu+A6MxrlQvY2ZPGpDuEC1E
FXhtOo+UxsKX1gF8plk/qgiqoSYf5wsAcIZmUEsAGZd8j6AnR7YvYBbF9ViUxQUfTdiHPxHRTcUb
sZfcr5MAF8JpgW79A6gihxTSzyP9O5RTQL+OUIEXXi+o3vBmLZQF+kWh8ZFnus5GWKT//DL3DuLO
eMgdvlcszPHcEF9a457lyGiWmksDgxWHzogwJpSPTjUXi2qUIVcjQb4/izTQKCVWBoLSyuNsZFCv
5FZLD37RGyzMndsbnEmeJ6FoF/uro+PhETTKJEd1kPTl2tYg1gU4+jGRfbSwJbvrY9HnY2da1jQv
X+StTZ7JyYfVETSWhoYVkZodC2G+gM80nkgqjwTtXOm0arM+04mtuGT9GTXLFmICFWtlCRfhdH8c
6y3rggyw7gtPtSFXMDeLPR9G9UHRfSX48j58Y8Lwd6dXubCt76uIm4NmD6Zu//n16Mj3UahQyCYH
JRfAo0abWfMYvDj6TxEeDqIv29Sjx4NCOjRZd9KSl6AR9X3KwvTOLWouJky5m8P8JdHkWeqWK7rH
R6f86B2W8xEEvYBrOjaqri5lfDY4unw+6YUWAsGDQ2ltWrCWxOF0fHTEy99OStUiSzvKu0vpHasB
gZ2Ft7mPXpYd+kzh2B2E5AXT/2NnrhhHu+qyaORrSu2aiewB9KAwLV6o14DoY6CJLadMTJ3dwJg/
xVTGEdvq31BrmPwITrrkCb/bGLmIB6TDNYKuT7DERcOr71tBm4qNnCnUT0zlGkKljSGpESyFrP2g
AZezwkNMxCCPLgYx9RMiltTUWvakubm+nHRXlNEHNajI+DZbzCt5trrOnADwvbWECxMK7YrQRxEC
LZVFOu0WwpY4bN9vq2H1CFUnWe3NNGfLuoIolcHDHnN6/HKaH6ASW6ca8EBlHH1SozPCI73yk/NW
Elvl+U1/m9ngrOhS/j1UVU7DfoMOa9RtvVPX7r9EUWWAXYUkoyu2jtMyMVJ0Xp5+XlOkejfFz7j8
ZwJufupe02UVIWojkLgsVJChnPLvOQm6euFil/kjBQMbSFHaSAFBt7QbHef0SNpzS1ZCDcnXNBM7
GXgg8oWfddsHl8LwnaISDbeZX4/hXI2AWu45CgY6Meex1oDbu5ml7G39LSxbgXzFkC6QKzMjfbH9
LU9wTiG2iLkRgYiJ98g60iXsB/xO4LtPWr8PdOl8B91jM9XIbx5J6cv9rcCu+knDAe4CKJCnA1a8
FflbkhrzuWYJD6SAAPsThcZmY4mbKJBLfIWHRSU5kPzLOKYpiKdzj92R7246OkWB/dTXBq7oQSfS
8t7DnPzzrHvOyCzYMJlf6ZaeMWhhwN0Ik9Me+7S6KwG8KvFFa2DKxNGEEykLzwZZ0NJM/407IhbS
jBFpX8QYqYks+kyZWCzBneXyfby9Typo6+8ajmszzVL4E9jTyR43rBwdoZ1ZYpbFiVFIFLSkwyYF
oj7bYShl+4wPkMVA7QaW3xccQ2HHgXg7wS8USr2qgt6g4sSGBDHKgCVAjbv+ZiUSdjbqywS5PGio
32q0+bGd+p4w/GI2hhqnErG5F48GYNTc8U1eBW2g+YeG5ypI225iqfwBGx8P/tTCpY2LmR9OTVPh
zNNz5S5zCltbtwZk3MkdMFk3TJkg2Hwb/y63gb1jU4YuXS9KL2trDQrRTUZTJQ6ZytMmFvAlsa1U
QlPleyyKoJkcyF/cFC9fPNJeWXqsqOQ+VpEA0BG/8gvtAEWvUCxrQGAPP9Y2jrQX9IgDhF3u4Dd1
esk+HqujDB9ei7G1nYjsgBmll/HloumGsSIdlxo+4K35EnBD5UqQqHATtl0z0Q2a1BK7YvVD9pAP
uxMC0QNnjcY7O7HO17xsH0rDtJ8N5G3qTtM1st4qPduotKAtomb/urv6hNNgPNK7U6M8ngDl73+L
eGwc3eQNAmo4vQbJpSD35znaygNJpGjqZNlolE7L0RKVayQjNbkAql0KqsmBKnDFjJYc8jzTiaHZ
0S356m319SjT/GCJiaxc65YccOCOXicrwHvTPPrjhDxZMzm5EFTPzVS4XTrpAU64VvNayoLVFjOe
SdXJxzIbe5NhazQzEYmEd4H6hA6XxUqnOaLKE+JI9rEmNKRraDE1kuqaJfc8zWCX2IjWtlRDyn+s
L8m29N7uLIDgnPSBTYIY1GICd8X24P86jQGTzuC3KilhcKmowf6Ld5ioN2HmnzLozCMWaKaRrck3
l0FpdLHMdgV7G73ellPtYK5+9nWc/g3sm7k1YkkjdG7J/Ey75HdzmIApAGbGQ8Umcl5HGQHlgR66
aVCcmOCHncp2Hppsj4C1pAQhYdeB5T6WB5wKZLmzJqQVkTt1pM6d1MhPsWGD82oimD7rBEKUM6Xu
yYBZzIpSuU63xF3618B/qErQxPRfT6+xk3v80oCJeVXcX6XaS55UmBKloUHld4x7X8QrqOp92qaq
68nbNRTxEGCMY/w3GfvhPQ3/xIBnFEFLY24tO2Gan7fpIQu7eOgDetQoitiiNob1bbOcQ/zB8KOR
7JJ/+ZVZuvvoTZkDEPnIh/wqp9U4zkeLORd9WDeCP/FxMv6YrTSb3Y0SQ0aeA2K7tnpr6uap2HLE
z7z27D57EZi7UxHumhK5UdSPvzloCu3LO/xoWTCpiU2Ulxc9lrQaJzdJI2khQmtc18Dm2W6YfCgf
qbkmAMZ12VpEDxfgs11jJpft9nN03P2/IHqS1tDq7uzNCPZQk0+XRkpj2SzE2Ig1pcw7AE3gRw08
61tf4i0HZsUouCvNlzNBHGrdONFWYnoJiYmMYIxnRJikjsrVIrwj8LX8YwIncIub3bkoEdvKMaDm
l7mfX6SuKR5QoSdghhENLLYtPBp5HurkZxHOpmkkj8gM8Ov8YARa2Njp+Z24yrG1ljaTD3xV79HE
DZw20DPVZPmsEpaWKqbgwM6PC+QXv+1jnxXAv/6pkhfH7WiLZ1rGLsNMXcM/ylI+PZ5PW/3qEnJK
hU2mCD1yrqlgZqry11CkQKcs8rLSshF3HLj891yKbt/IhgzrGSow3C8OdXqox7oCvMBuh14IKnxw
uyA2igVjt2h6yjKfFeb01c4fARf+Z4A7C527WwzvTHdywjAsSRV7NW/nMIIDSN4C2DG3i91WETSo
rw8TW9EW2muIBGmlDRGbLnwXVLqFy+F376UPdp7StVaA4KoLuEVHXAmu9t4sQRU1hVSZL4+yO5JZ
J2EWZwTvj1k0XY7bMGBymGeOx1+gP2a9DJiR0a/u1EE2hCXj1/Lf+Nf1N/imwJvdqK665M6Fgvl3
8kEvys39o2ZoxFyCxNTYDPLD3RcnuP25DIJWJaLguD6vyRu/mo/snE5aeqVPE/+t9HT7tRyNT5Af
CMW0Iv2c1IwHQTG48HdmwNSzK0IuwUQcEmyn0IxgqS6XzVqJZcpCV3Nwak0y6v0kTXf5byM76vnA
bX5NpXvsqGpaN5LSGq5D4g5lAC/3euUmsnMnRkskyOj5AiaFbepfL/dYfX2f40lAkDBcxywiMOSS
1+Un6PWXeXjV+VsC1Wcih/i/9JE6ukCCqwL6Laxz1CA5ps7iG/WbcBkQiOTgx4LCojiM7jJ/mfkk
5ZtaIi4iBhUZ7MBT5CQmJPP1kyrCc/WYONZUSXXRff9Etzzw9muN4Se7WXN3pQI0mwPwJJMTNA4b
saOrJSWtnrGrq/hpcxx8qfBiv4RF8eIlaUE6Dts7mIKSW1EPk/0sKqpMGteLZGsQtBLYVLXzAkE8
V2wle1XS2CqQjjGRR1Y9rwyGqPZX33VK/URN4KQEaoDEfWB+UgZGAJGD7+G4909rEfe/DiQ5G+bt
04xA1Z7mndmN21QemK2A5h1+otpVzVgk6h5o61tTj6qFuDUSXKWr94mbuCpYkaFvKi6YZmbKfRgY
qm6GVJED/pBwqFfuz/4OdnqE7jHqgNjBZrX2J9t8IjfvbZ296sgZtz4kvV0c79wMoE3Tib1YnmnD
95mUNXe1G5CFt0qOzQx/g0Atot7xJoTQaPzesBbWohac/1y1R3lzQaPkqyeAXdEzELqGv7VQ9FtU
LTY+np0Ky++OnCxNBEwMRedzC2y4eWnkP3/LC/9b1jMvdPWNB4mp9sxXlssaK8rteYX7dErw9u8W
AQGCSSvsuzoZR5PFYhMUbcDBuJ0UEsjKvEdGX0OTPXfRU1Pv8hmeJP2ndLk7rj9Mnt2qiVeTA68Z
QX7ddYprnGafZREKddUnKwpJiPTbYY4hgRMU0NHp40tJ6eLRbSr6XB9/Ame1TxfsfxH9grjVPhVA
0kVhLH0uP0Wzb/vRBC4Ok9k79Lse4kqgk1IG03cOTNyIHo734cxzoRA+199Lemdct0SAaaab+s9k
FO9sztQlBIcGsr30+gNlIIcVtDlcaD6ClHdZ2j9YW9VjR/1PwMnV/4MfD/xqPqftgDo1gLQwbeYL
2xjEucXbdlSWReSrjulClJ+lvWoFBsqn8VZ3AcPWHxzFFjhsS0nxdOPP8Xq65DZYtJQGRiX8UlBA
zoYRIYTu3peBsOgBGG4S8EbVuXXO8ajMjtclAZz/zkAzuqDo5Mg78PLiV+I8IkOoGnA6ldCYhnOn
wPwI6gJ8+5ZcnvgF+mNLXtTDo+nZzQk3hy7G6ms6ACnLu7etaeYfgwfKm2Qru0I8K4UV6sFPq0/U
lVCNRLtkVjjBWsUHxMjvCxseAZXtEoYW2OnmMKelh2BdnSkKWD4zyslPIrDZUprIQtXBW5Jt/AtP
vMXLm0Q9uQgGVUbuiJiip2lLPK/w7CGrREq0T6caAX0TOyQNwZxX9qkSCTvCAZa5N2+zarH7RJ62
iXMDXrqswQfA8j93XG+P5sKU3z0lVNmAbu/IP/YMYTXgGACM7La/j0rwG9r0RBD/UYDfLPNy3pVE
S7KW0vkMTE7HdAXyLaLPZQtz+2LncpqaqiOtPMQ7O/BZrJ2hOnDZ6MOwZ65eoonvpI4vT3gD9Rf0
X2TcGMMt6GUPZFuR4EZ7dyhSoNvVs8MipUUKRxHTFupvLeq3mZ3OZR0bB0t4PJCSQYDBmbjm9vNt
n1JoSL1QUeXm0OiSy6i8+xZbGRYHznkAYwgm0EJUe7ZknErs7LV46dI/Q+S3xi45lTHFSprMcJu7
RTDD4Q8u2Huoo7664NtUuiVTwcaHcATX/VukOQ848UsGUrskXJBrZSa8MHBzm2VLrFoMwIv/G1r9
II9Rfk0b3oI4YpmUggDLm7gFTstcd2Jmo/byEo8/dMTP2BoO5UAH2VGPCVovU5c8rf38tSXLPU2S
Svf6IWXfK7o2oOLuZv+6C7zVwRf9O6Z7MSQ8lw6NGGRZtjb+neiMecqoLk1LnL/D436/hSzp+O7n
KJ1PUlGT48dJONCqrHFjZBhOTgGb2/+0kNVRJsN/Kctjjxrq3AnhLkuqTT0Z33Csgl7hsjy/R0ZY
BOm2N44LvVm57kmX54AUjlhy3MXtyA2OIaZ5JNjVmdkQiSp3Sufcdjp6XnhvdSTMKI9oFZsvgEXO
MKj8F2Brk36S3IX+U3cWqc4q+NjBvfSiPS437VdxhtHWrb02NCJVqdYf9FYLY5p01pOrP67NuzYo
HtX7FiHHy0JSgcPYJ4s+uVLXAxTa8IsbNzs1YsIwurWaOczCX+xu+LazyAbvQIqp0KPPMh8VSQHd
hfIjC7Qg/RLt4vJ8x/DSGFk8OD5srPp2OK+EsFZgNCaRMAOu05hrEfRTJqmO2kPXnNsRv0qG9HE8
8nmcc1q5G6giCoH8jHsO5HGkfLhWoSz8yziMzn5g41e84peXm4XYU9uOUbgzzT1TwFVrJCyfOnr9
X2OoN/0Msgy7140bfArH2Iz6Lsnn9MdHq1ZG/1RCi+vn+M5XIso9ZZNOxZyQ79aJIhkbQ2FknSMq
+RmTgwEXUw9mvG1OPRDqAcVrfY7RK46wjOqJL77N2/ATRXES2Ft0BnohxLQk/TybF7vw0NXXvUQr
Q2WYCaRt2gWcvp3WFklo7oBQN8kkARexbRfhYoXKK25absIhEM/eW7nNTFyfcTtETtTu3OaRSFFn
JGCR/Hj0bxSE9tIOjlVDEV5nyel9tejlAvydPO+VnV21mtM7TzS5zDLpnltHQP5GOulqSmFLPLpE
hS3w+9T413hKHzaLf0ugNQ08KyYy81MWlWQJNSyAf5QCdBMXhFT86Xx3aBCpSV0CPuecE0gsje4H
UIGzx7xDNjlC0fi0ZW8n1KIbMeAkxmJVXfgPKZIB+ITKFOnqwA1MFqKVCEk/ekU2Fy9HcUz5S484
+S16avVcmOY/mwulG6dtY9P7zYeAZrma7FxRlYsmB7aM+t5epGcWG7FhCbQXJcYQhh7gaQh0vPlx
+tNkQdrB8b897+sEcs4Kh1TpsBrW3XN5Exv4BWKqVBpIvkFBpmRKiMywMD5Zx9tS3GmRbJ0Leuoq
ezFI+Y1dwcvzm53/M9wSrnxQpJVLwoqNdD6gN1FBKBBBcnExuY58RFrVlVWF2z4r3NwxrMsMwwKk
VIicts8VxPuP9b20usYe8Nx7at4niuzQyK2BIvCoFimz4yXd35G1z2GMd4hQltvi1KySEanVtKbU
rBF8cn4AtWkQU7RUGb+nkvY83Pd5lWb/1Ua2BRWfjiI1ccExAhFL92qAF/4RO5LryK7YdZ1Q4rYC
TBvmNvx8hEB+DaW98ltGfBsuI376jmYg0235uQZd7KbQg8XY5Ko/IzO0Zzp4rvuJLAo7oP76nKHx
Wjl1Y10muEdrxGUzwrF65kyttoDyWl3uZOxfCDdmDFUfEKVyWJ/mnlGiqBQYkKTe2k9MyfmllpP0
LpzphRbMxcDWM2cgNTSgEi7Pd1Cb32r1xYExdaaVLnTF54RCXBFXu2paDSfb9S1TXDSHy495TSPF
6j8rQ6vZ5v5C6biTXf6p2RXT/tc2QRsay5KYpDd/c5vEfCUVkd06TP4KLywVJDDBOr9LZ9Ea8Hsy
owaDIVIboENYrlNaxDRwQKilJUDn3Ly7En95OEU7RYnXX7O+qtSYEtcXeySXfOdOr/Qsa6l7bFVQ
AbAW+RdkTCWGKtwZfaCDgks4G6pp9/mjVaC4nUgTVAmh7835qKUxB77djIaCwAD5lLWxlYimFK0V
iGUWuoRfkv65JuuARMMJhwlcQ1qfIqJsb0laJpAng1tmDhk3Y/YKym7TYti9MsxiUUnfD8i8ouVl
i7YApNWUgSQkjb/SoRPPx4MDxwtx0YmrzSnSXo/1dKBybmhFaByYtULMkLzHmZP75ZjRePWhS+3u
elblunk0a5cGtuoaqm2D7nPNcThuVC6ZuypCJhXN9jDAhrE1GV6XqtEi81taREDldZmjhMvD2egT
v37xZt69grGAPC7ktsBdr9QrKLyyGUFAEfrchFsZSrORLR68cPrOunNSpFP40arxZiHhoyUUk58Z
dw2tzrfw50J2kmYSVKValYZNRdRCeTDs+AKi0+JPKb2nHa5RaWyGVeV/THo/ncuriRho1uwW3VIM
i7bx63GAf6hq+KBiGH0XEHWA7CY2kUOtlgjBoVU/eiDm3sDlxsBGvMO7hmoYpmOkot81Nxl45Muq
1kKiialBc/LhRIEIxbsHwZMWWGL+E+i+B94c0uDYyrS3+a7ziUC61cTXN4sZFAR6T+Sf6W8xiQqE
eAoV7IR4xheYMduvDeifLGob653KeqWzmnMyNXIdGGWa11pPN4zIfFel5CjQyHevU7xFBdRLlm50
8IiyOL/5gE9Tm8pxT2+mLvfr+0Nh6019dtKQ2JgD0r49sZlX3exDspud3ort3UxuOviJ5H4hnO9L
9kC+/7bzXqtR6dt8/i9YXUwCIZNKGnMTTozrkYDknyIi16g23j69/uCHnNdXt2WaDr0FZOBApx6k
49B2Dv4xTdGgsZ0Qp9SqVC9Wk0t6EMoyfczLgrB5D/2qYSpA1nOMKBycMoSTjPVTRD9hVc0ZnlWy
Lskv8/UKemUJSmAQ4w3AqikXT5Bms3VgGa2EQQvQn+FHvjoWWc24NTtqZEXYj0t9DgSXhrvOQusD
gYiwM15DB+mdkYJrmoU13UuF06C1jxA8F1xFF6MiqFINO2z2xF97JH4CoZX8zQchr72Nf8h9LARe
vRKcQmpNQD+CIgahfZ8HTYmmKAzUgXYNZEojB7g9rcRHvBC1SGtBxVI8UlA3hLC9Q1sM0f2Jwinx
+yQMj5fGKTUMgim6Olb0v7cbLuyHxdo158IQZAYsSC0yfElRYuhF6hIM2PctA9ACuKMqRdhm+5nW
6BzLS3dcRHqx7w+MrEBGUZnGBHFV8FNMrv6EpIJBBqVZwDlqpoFQqoJMUGmhamTtIZUhoIMRlnRy
IvuTpIvq/KqCPOhFA8PVHaGSRiKCWG67yQwAu0cy45wsDPkg5S+X6BAtA4sTLoqmkXFwMD0vuyjd
7V7V6oi6MrzaZYDfIL6DNw6iGQSTE/090jUpE4Hv1YdoVjzQk/lUu9PlsMUbeJVCDKyVAcW+Yil/
Eo0cMhg0QdlZt8cwbYNJENxsKKZ76n9ZD2UeHp8Riy1WfvdKEF6EMn8D7zWnRLf8/3olJe7swPNs
h0zmcg3j2ChUw3uHMz+8hp67F9RyLQzY5wxAZ1u5yUmL0a01YePQUNZhFyi7IgabUt03S5UVuBD5
kmfdh5lzb7/lmbJfgEj10NLfeCF1ZA0H/iYIrlFz5+niAQhog3e5nJJZ9XLs6jtQPdBda/gSkdn0
zlPK1d1VCT4SLQmmDElee69sBwm1LvXZOgPJyofpaT5tRZt+pOlx3D1h4uZKgHaFQgCt8v84q6iC
QOLvSrdrOf85yvvCpZj7e/Rwfwihr8h3y4b1YkSAw7hG2iBFGh9f0leoB/sqft95SyZ8qAwnPuy8
6eBUCvWgRR9DAmdd5SsnAYXtzZdlEUBgZFjUEIauKJFdCzeJnV1UJudYwFewU5/hEPXNLzhbkJOo
U4UBtj8YvzDCWLdkmtXq2gbJDWsxBqHLppVlQsLq/O+nGF2twLkr3JdaLegOX9SQhNksa3w42VyB
GS9xPEQVGgqZZ6KwoFaaR5+tomnboWfIwSjyclE/iZZiDFWotZsiOGlcccKAvK31rF+9mzLiK3pa
jjgg96JTo40DooCbfI/sPBShsewidlaNnxduVX3RZPLeTmTiwQBmPCrtRhlnB1omGUTGwOzwcjBx
ePnVxRfa0OmCaJ0r42MJ54zBUX3leDGFq5dzTI241V/LD3SDQDF1OggkRXc2S/o/9G/wjQgGBFOg
6QPcnJm38a7RVwu28xUdZru3Gc0H4CggKFPO3ywWWmhHYyUM3DiUiptAgdjkLjSQ+5iZB0V5OLCI
EoeL+hWfZp0spSQ9Fuv3B/5hq1UvFy2PuCJHVBluvs/mq5JOL0NXKltbh2g0qJ/o5NPzkgqQp4Hv
QFFzTJeV2uDdkIbYMJY2WPZuq/gMh8v/3VFmM+DjwALfy3Wz9VIO3aVMHYAB4P4CCxR1tulWpzrQ
idEvOaO0uPKSyLIqMcqzLf7G75rKbD8MdDHXVYjEnfASNbjd8tXJcMibDifmO+u46xp69iqkw+V3
k0kwVAMmud770mmoHiZiPJZTM2rD78F+C4xI/1BDJDI40w25yOdEdUKFVp4KOCJNj3OS37wNNlZ9
9Fae6ndU2jxxwnk2o6wwVbGw5fbE7AV2TB3EpTLYRFi2PGwJRzKzKaMuwtb0Sv8DAWJlRiG7TDpM
DWplesCPm1Qm5H7s3qAHKy2JyFfwARi4DI6w+XtFT3NRLlVWIjakBZwGrnJqUJhkjtIg5CAa+CGa
F0ugKVWXmO+ra0sdAlQcderfh1mhE/VMJhZqZYbqP/CXPBgJILJq2nA3Vih4UvEnxWPoLeg+C6cb
B7OJurXzng/ayk3UW+aC4d7S5OTNJgAMXDqzQWHXqgE6nLKTiIaNEat4YJ4Y2ZaNWTyj+CrqLWbv
J6shNHtli+zQMvg1mnO/OKg9UuJqP4FZntOsgHxpYMOxPh1sACBHS4rAI5QbjjJxTjFelyiVL8iJ
R1I1NldMabRrFH2dU/rHlSGoQeXuBaPmrTVuMfIBOGpEe+QaYVJqF08+fnAr+3mvVifbg2kYtLUL
VeZT3AgbmTvR6Bo3+E8UQZK/Yb3p01wjbF0nbVUCaOpZoshYHuyKxlHl8qOcjCPEMVMQ/Zpp7kRk
jVM7oX4F/EKiS8EvlXJ3P73Xu+PVwK1Pl6/QKT9HW62pBDgJQr7D/bwBAE0dNxoP4aVOd/FrIfXa
avGRhJXGCA0uUuIRo9nqe5WyyOB1vM8dc4izTczH4dGylMXM3VnfeCPD8IONIaen6QAa631t048C
6eLmP/8Mzjc1YfBZ7wF7EJ1lxHeO3ZHJ1el1KFjHahBsfiCKA9UL87jAx83xrWf28Wvsra0mbN7T
7bGJdkiVXZOGQmE09EIRBzB32hkjYj6n9WGXJKsVbSto6RiM4v4Qarq3pms6KpZLLNi96CZZLj06
ugNT9yjIKIAmM2pSsJBIFhjs4/RCoYbUcJrcVGEpPuLlbZ33p0QbnItSKTa24FmlyLak2Xyb0ZrM
qUjSajSdFVjN1lrjjrIxonzI/lgAhXyX6COcoKGjXkyRTrmmnoBqzKUgcRhiUYUZzwj73aFvNil2
mQSUxK167VL4dmgPSSELg3nFNLFf8kS6+Dz4xlUCiEfdsLsb8ur1XR7pgYiiozM6VWeCuwqpvcxI
HHsEt7+WgQ748sJLve6okzTwWaOdQI9R6Y+wDsb4YzhnDcbW6dGQRStMCtA2AD8Twez0FUSxygV2
mr5yT9O9iyc/Q4U6OGp9gf3XmWKTzpKpRFW4is4jPY+M2VNxxjTo4CjS5y+3uRhnCaKD6+vlSFZF
RvIo5/eCjxxqObeTxPMdt4NKnVPH+1rqYeN2qwFthQbzGyKIxLLkHxTgBHLmev/70LfPIVXGdWIt
K6jWzOObrXkRPY2eK1VkrbErp6E2YV4Cx5d2/RXgWdzh32uYztiqIdgOFguO9ANF4/FvKg4/TO9X
m4GKjz35YxYlbxA1OR49FHQVxMsQ49C03Ga7l7aOaWu0de8huMOPDoVH2AZFVau1AUF9YHJfXaUE
h8BKJetrrVQrkxGqsdcQJLxR/3xnCUhKqJ/mRJzXUr4LZtlOzP9o+lVLOy5pUlx6bJEddk3PEaKI
aYrlL7X55i8ZR8mZtLvZEhTOLNgo6mbjviBv364PezZyo7jaVOGGTsiXkwh6outgfxUgEpLSeJfh
PiIaD2qVvZhN9VWoSRvdRMjca2UFnOWVEdOGlLO/1BA/wS7N0JecfCmvTHUjCuYBfvFWrVcuGGZv
JypG/fnBQB0QpDl+JpgAx9MopjjxADYho4PSw7uhnJ4zBstFDs+EZWJ7s26VvOf5VDPSP9ikOmfw
NTWqnXRguz+68M86pUnEP62AyqPcN14pZpRDnCan4NkZ9BLyvlx0ANm+UlKfX1FE/gfA7ASujKDS
8FiwEA72ZYFV2L9t7HxswYtwOJRhmDbZJhWbdkiVE3HX4wgV815M2XWH11OZ2CTrfYWzp+zHulds
f73PJX9zjK/c57LCI1MCww+7Yd0J13/gEX2ikeW5NrvuNHhfReaHJR7T5c0gq8PoeGzzijjdYm93
2/oTG/jf3HGF8b4bMnj0jyyeVodvk/wtrrYFN8ttCHqrJ8jMx7xYgUrwLg1nm1N0aQDGEDWsb1wP
wt6MmwU4+dF0HW9+RUtmcHYXcsB3Zqiu9fvMXNvrn7Nq/BOEAFvKWwruOM/j65xUMc2r5YDlS1nd
duKkesYXbfoKZyFfsdqniCwi9Ag/pwDdGsh9Clp35B+jzv4Hgdz37yUZPSceN2o7IFi851+hcBuy
WmB6e+sUbOYZ6CQCIihWbQ7QJnkx1Z/zC0Sy1DhvPoELZMfsYSQxDH4ZsBvT0gCZNRV3QuRIifWG
5/j3v/17QxldGlZuuGof6ZvhkqvqUtxoPIqEnUITquVCzSie9pd8mby0dmpLf2Cljxh8HC2Epxy7
ZSoPInhueAXF9PgDxL7vEzg/GIu1xMppkXmSYq/qlg9P4d+t6SOJzzm+0R2X6T6NAoBCiwmQ4JOt
bOWeS+RbFMdRvvmH3WVkBjW7StrmDn7zb1oamzqUgiGjWDU5ES5HR6zxIQ3O+5ZbGNJi06nLuTvI
UbvmGhaB+ISuZflWUhCPjVkk5gPFaYLho5vzFHJbJoMiexxaxmW+tLiMuAGBb47O+F/2pCQk9rv1
qRDzUtcayNwCKYXnoeQqvkxONztGr4B4d/wvSeGxafK+RkVhjwz0d9vMnondVMYEqBMYCayel3+Q
PKoQ0aVF6Z+W567V6xWL28qLSzWvcFkYAXn58gcG0i5e1gBBm+W1y/MHNHsjLbncoosZS6ME8fy2
c0uSclOxdde7YE8lx0RFY6BJJc/ThLNHvXac4RTB4J/KBSXoFkuX3e/rlz0TPAld/V8dPyQetrG1
RGgMuVg5gVJP61/4Ckgv2j9MmLb3zY42faHXGvswPZ/JFH85G5936ummu6E2ACipyISqpLJ5KhLD
wbCXVeYOgLiZgbE1L1slModSq3nTqM5qQNPzK2SBcIUds+CsfYoMQcPqmcCVGxEHq6ImmnpwWidw
6uzFGu8ofH+ha1iMFtaKA8mZNdEaMEOhA/L65KSeqlD5mn1aeEE3El6KERiWkk6Pv6a5cpFL2Z95
tnnJG5dk792oyE/J8AG1ioWCHFPgxsHn09QMKAe/jDB5UodgwX79OPOCY81aGEMZZl/U6Qdww1L4
YlkrnVdCgjPPR0IDPPHupHk7LaB5L6dDjxfW/SkdwgSJqiAP5X+mwi6v1wzTnV/jjCkDyRRj4IW+
oBOoJZLFBknHJR9OYTjZZSe7aHeGqEq1JN1gjz2J/AX3BtCLi7Tz6zESxKVH97zUXoreHEvzaIOy
cwXd/hZsyGJMeGfSisHePM0JfFDrgpjCVTQBWPC3KZgwdKs5FbNkJA4NVU2PwmBuRUO0lg5HxZld
JuLMHVTGcJR7Ny5/ARJvyC0+rFmlUklSR1EsSwxmtNTT5ZS5H4LvHNEB9BpZXJJeZJpSiOIVlwKa
XyMAqOWfCerXWfNOQ3zTlpyVT2YICBkQV4dP5SOBB3tJq2s7eLjOPWPWL7B8kKSoI5AGx+h13aqu
jr6b1ZghDOCJ+z4H9B/4auQxSinqidrqFsEYAU/fIuFlZOu6m4iLaFXvs+0Z1i+Co7ISjjEto4Ic
hIzRcJor5GO4OrpZhVHJ3OBWMoEyxKDUfflDi3vJ1xcTNkyZ2eGgjuV8iHAJm9Jbfd/1smB7xj++
mm2/LsZqjambuB00n4GbRbSz5hUF0XRWB6ppg4lif/DFaf7E1nu1vwgmwn0wzeuu0jtQoBzCA0Xl
Jim420bAwJXZcWz4tgo4+4AHrXVmJ0cOCBJy8nyg93R6VBBZuZBsrqujwYySftyPhFcegVnSS9JH
afH4Jrrh5TnYLGoTmzVwvnZ6P/fKvg16Evn2yzM6NRGtbIyZf5pWdR7kWirTAw/CkTPXzPK9LLNW
oLwm3PTqFSPEa5G7uvzKqaNrR1SN1aazYFMDq9jtNYDtvXypZI31lsUrJ6nhkY7UtsdU+TKhyDcA
khoF2jVDjLm2aF8Y4z+mCllgXDTTnqoUXPtF6mLBcw9mXtY8dSCDwoYgq6xMCQrtCLaK0x/MYeOn
Pdv4T3FyalxlM0HC0RNWuOPsjHJMCF/yfxegRCO7vCIVpgd0uSuuw3Fo1yuX2v3eDLTeXQ758aCg
AZ4WOMyrr5z42K8jueDQ1XDTopKqVFA/DBTvvLPiFNbJfKkueFT7FG/VJ9X12bmJAQT47kYcNGdQ
BF8ckmwmKdfpT354t/AKYMyYni9hOCqQVtTXigr1d0GEIoTcP45X96Q/3Amb/ClHFkgOnV/aQuFF
cV2kjECgHjOpkaGJPScscnB7Tx1vbE2dnlPzOcXp49QflwFT5Hh2tKt1c2t27380SJMqXl/CPblX
JYJ+50vlQhe62+z4wYW4t1I8ekV196Q6B+A++8S2GbOXNIg2WK+qfSw/YNucpJnccP9lbS+lDhY/
62FM6wJU1t8fgUGWA0V3K0z3dyHCVdzHqHGKFxavYFThWg/opMhHgNBHA1R+NaeUc9IylfJ80Es0
ZY5VXlDCjUscGfu9+AS7QdQObRlGh7ieXBm+1AYzMpmMgtZ7A+9UQi1+4U8r1KKUTnoS8QyR57uz
1Xhaf0Ht50+Gbwh7g3M50teXGU8ha45D920S/Q450hDwpQfCtQprL25o2tfehAZ+4jyZiNAKrkA0
f5jo4R/lzGlNGhiFrGFPae8K25YZEfLZ/v9KrGafiH9oDaqBWQh4e41KFCoeBioaGhBaES5jCtk9
pCdx0s2yckvRKOVhLJ4Smpt8uFCIjrjzUCf/wCvqwdOdTEkAaQ+YJxGvJEUeBXHrUrra3qzilxHE
g3NAiD0fhnoCtTihgx855toKojp7KoL0IZ5DeDAizyLtD4KOMXjPUhFyBlU+RRv6rZ0TkvQfS0T6
Hrq+aVLydhWEqbgCGr5TJj0NMKC7umnM3so7W0p72iGkRGVMtrneAVGtwQCjhvMnK2wY///Z27b7
j0IC0JkYM7imUbRY5/kUm194dgDnZL2RhkuRP2zJ5DTeE6nRWdBv8T1d0nBXvZXfSRKfJUNlB/rO
yklPQ83s0GKjCd+ReZzskF2+jRtfz9aSYQ+EwjXx+aM6BizMBAwbUJN5navehcTxGXN3E90OOTSI
ZaHOoakSJ7uReFEsPTpvmVWYwrU7W8xXydUZAqGaJi6SYTcN7aCxQpMBil1C1IW9hmrCoEquaRDv
py/jzNpoJrRZVEtGOPxFiy67JK0LWLeV5Npr5dUY4CHq8EM0E6K5L7ZaCTulpJSFX7pfWn+u1Lt9
ULDEz4B92Z4WyhDDURcFrD7doqaFvcfjE9egpKggUGfuwD2fYpsBPvxyLy1ACPxatpA/Zmr5YUrA
fp1e+H8EVFcTo0awbJPVtbEwc24iHGiL/U7oILLhKeUawexFeF/uBMiz1F/TqERLEPXDWUCaTPtk
ni83VxtzJbGl0eYxh2xDBiU7HAau52wn9I0cldpX5dJ8iOul6WvLCNiF/SdTQkh2bXhf1vj/fdlD
VpHTFK7vNa1FEC+m78xdEffoR0ukMZigt85F+tigaDTfkrxrpdIjnF7C07f7T1iU8o6+q8/yX5ct
U3FCibX1h3YRdBuI2mM0XjTzc0suEEZ/LuCW0dULUFoJib4AJM8HFoE3HpxmXUDcUPVS/VgdA4Fk
npjBGNTjux/yh8axyRF6myQ8eazBIQbpABKrQ92M8lAfDyOXTfDNXIIijfwoA3TQRO0mnDqPKY7t
GKkvOCk5rcSo2G06KOeocOVA20gWq/jrijQKpZ46ciqT5uQL+s4UHmDhbGExK9Iy6u9nWKwaBI3k
xb9vmPsD3nKyhhqDibpZ9ao/tqWbbiHPzH0PRTS3Xzbbn9eNOTiWkydgw4jaXhoa1qBkG4MTFXBe
o4f/riBFTyL4vvKphKfnEs6raw/ePcRBfgy/3EoQaSePu6KpzcrVyU9kdvgW8KKY82CfW22AH4Tt
4ksWSBZs5PGQzyBApJpS5YNk/67AepHFLlIsXJP2QLMD50c7WGUMX59N7ARmvgqz5SQ+0NNL8aPz
fDSDeYYmkKhnnXCkKQU+mZgvADfSEnOWh6uuI/oio4Xc0GcoqG41RNrE6LSYATxNbyoIQ3dUpwup
6WK9U0eLKbVufcQjjHopoH+OZT6CG+g2pA+FqqFRc8jwvBanhO43JVsx8t9OjwFPZbhXePo3tGoa
CsmYuhjqCHpn40zy9xKHesg0pEu2MiYdJ6bJJAFcCnBsdft6nPGpfacqTP+r2gLw3fij96GiI+L7
N/SMuTZxkD/PL1hJ9Xxa+o/vc+XPPX7fZKwz116OlOKXNoIgRPqxBvXADSQ//QwrMl5mK/GIWrWt
WZ9jHC1+Z21Jdkmn0UXoYWTp1ZXiyxmnQZHmQJucUWMcGZxsbAU9iY5hrIkExeCYmtHTy5s0fh/D
E4HXCxnMnaNuUUBQ+QWeam2xjLcKDzYFMdpnnbanwxcugPAjnzXbv5zfJQQEKlcXt5zKW4DvRiF8
vluGYFn+XAi0IjiS1nbp5mk2oUMCu/JvJ5niMmEw2OQgRtIHNEdJJi7l8rminqIEV0oRkUseFbjA
neIDNESNeU2wWNJm+wUGGBiPlMt7+EXouC57TusRZmSHU3ru/jbMaxYH8wCdZhRo/5TF6/L9ilvS
F41AJw+qmHk3fpkq1XiqcYBrL7v+ChUUo0NBIS/MmqksokhvVCyT+fXmx2nILW0zfQMkDp7Y7368
CFLm1phGkrRSiatu8pGN20OBZ3tv06yGTmH/IqmNTBJm0oo3G5Jfrl2GEUZvA2WWo2w5qbLc1YLA
pu8w3pQArMOgvxf0o3Zm9YHG7CgcCkeRShm92pXzlXvrPUq6tYRSiVgDfQsyT6LQwiHzQwMrsK64
xug2RcFn+w7SDT5rUG+mWUSozJmdEI3T3VmTJUq9PgMcjn83CMuqFozTIkn7q+gxK2mp1zig/fQZ
DmTQ4Gr4fC4ObYuLvrFA7mFcG6eX+oHTue/Fgq6rr0H12147aaSV8B2VV1GzSuEvvEIBEls3/RSA
1nT9uDOl+tfDv3d9YVmXToJFUqTMkRUTLFdRIlva+djZdi+zryLcW9Zq2JzJM+sSPQt0vOlbak7J
Pv4qJpfG69v/DAcsWvJOHeVCLQ7A2m5NR/bRN0fw2bajB8ZO4x+/O5cMrgJtT7pOsDI4PRPGBIE9
IcKCCQOH8icMkYFTo9khzxhOa8ht+yyjWRS2SjTgH87Pxqtpwj/71+A8JU+/GWxav6sTUdHl7gwt
mGCNsA7t6/Cbz2yC/EA2A1vHNsDtooHAi/BpZzBPmzlQDjdeNUhH3b1IvepHWC/xrW6Q9BAHsjHU
ECBmnLAiqsAIPPWYly9UfKN/9GVexmivICu1BPiLbbQQmrC5BtMhx4c96Y5Nvzgxr5qKnxzPigZy
GaGVxGXtm+8EBgHTwMxmYqxcRaTsNYRAQ9nFQmlIM1Pdpv6Nl8k/vF72rTu/XWjmhqFX4otVhUSS
u8Z7on5+qIEGXHsuQH8kx/mznK7KCIRTH2WW9yFXct3DZdR9lX0ooqdrKIQJ5kRQVbS/dKEz1aXv
bhGM8Azdp5Os0VnYVC5sXcy4jI+UQyvnz7zJnJXihwi2w4i3vAe6ZFUdR9BK5Cgy0CAM/M3GsR/q
9vfL3mvuC8Z9j6JmOQ8757XoDH0yotfOwb7+sIahIHZvauG1wfskwT4AE9XBmQD7CBTJ5Og+PzzL
LnczgpLRdM4ShBwzVBDAsBey3GdPzetiZXhBAhBJyw3fdTZyenGKHqe3xb82TAIzZ6X2PUIv2Tjb
DZhWHPsxQSuqOL5fndSyeXoWR/l4S6SLiK3Z1G3fc3qdvumZgHpLGfainzEchIK8NCbIAUU0PT8x
/JrosfA7fytilVeJloDjNhiIsCNBKZTVpV0Cy8nEegtjStMoK2wXuXFLBKd8t8QPnd360GHfjYdG
R60RO6jzoEw379i7Yuag87CF3XqDcsmIJx7OqmsYd7VKphfIYAKjEtFX13wPyd7dLgeeXUaHvF6q
ChaC4x0Tw+3qdoQsP0zDFFmmm0Q6TPn6zpbD6ykliojPDwBWxjrxUyDWqGuX7iEfMWG2B9GkhfFC
SFpqZJamd40iO3DX5nd5JixA6cbC1eVl/CtcBPBuMOUgNrL1YZnFpnHn0G3YoSG0T/wBy0bRwbg2
bjnrOt/tLh01F/VU82R06aRJtby8Hkg1MlwuLGurnOnZX+KkoLuEHOms5VoJbyMTr4J1jz8SjBfQ
a1NuVYtVVh9pu9vWg2VcHyq7FXS0wtnEcpifY2eFTokabMt7tzJ9MvF6rvb0MKhNRX1oLU8qHJVf
ASMpDBTJMZDwCtbFiqrijqiVemKw38jXhz6NINIfvjA8VHIqGH8XYScFV8eaTU67Xq6JFyE8sEPO
bq7Aw67u/wYM831tCkoXWBvnWnBgq3C4dYV3ChKHofKgv0KJj0nlXNGPnnhLPIJPxhcL8aJcWGgb
tJJNWDb7m44QwpZflnvzbV5kbYtG4c0LjsKSXssOfamJANfMfMFzSLfpSyRipCtHbK7yvF6GMRE4
yDUYo7ll2FHxDxPBfFVKIUQH/dOZvTWPN0uESapUESrA4B5h03Sp1x1C8lejUe1b9P9VqxamAOt/
ACJxNVeW+iOU7XIEVsdR7Y3f0lztl02rSmTk6B+oD6ByUc4/VPBUYJJxICa5YAzPDd+loCiXn25s
H8429O7Sm1iYD4iQs8z7x33Ab+Vv7MPWmYm6BeKoO6BNQQ8DUurnf4YsQv2uZJQ4HkTJmKb+hHO4
eTSTc8VoH6mmuP1CWT2NgrLKDnLONqy1aRELdFEmSUWYJXf1p3yETI8uecCMYWFtXhOaOxWerEC2
EpOe8lLM3rpEedA1H/WqGrlRxnHknMq+nzDczI8RHRtAFgDE4gvjqsRXDV0R0vmLrc2UyHBzsndJ
UhJFRExbIXIaO5KiK1vo3+MD/aGCl77ADAiELfEyzUsxYLU7VPZu1AcG4aOO7RmiYiePaBj1lv6i
rB5Hu74GjtaJew3AFO4HNLqSNXQ3TooGQdH+MdrkSOubJ+cJjRA6x3ySxg7iPevcZ3ysEtqLLBCI
3SsOg6Ztl85kKrKFQ61jNVJCfCqdGiPfP2jtRSsTVk9Bu4z9HH65e9P95ZxqoetshiDESMcRDhxn
FCDqj3RrhkBj/BYal5wtQeVBPPEcNpZmH11E3Vq+yKBdxT+LOFcIsz6c5BDhsscJwYVAjl2ss42R
ynvMKISdmPX7iASwcO/AR/9PbWSuINjJ4PXVHFyKQ6iZQlW3Y3LudRYkr059ZQCWztWTz3p1tLLj
N27cwQec0p1ptO/aq7hv8/k8hm9g/q6JreUyzOnw5mFbuv+FJsKwdYeexwQG74pZYXF8C+iwqlIx
RVkOhk9nAgFc0rB1xZJIgorEfgk+44RtgKSSlgpmgWeOlcLq71XncNCyzkyKnlCmlzhqYxF9+6Mf
7Hr6rpakXMPFAIjpQLDPB1JVLRHNndaUI0cpPCalS8jv5fAEtWDaCHuy6b9oWB35csyIBEgXPV6L
RRQEzVVUZ2HJJVY2SXVQFgWfT5UYbeS7JWEBTvt+Ec8P86VtYT/5tuwy1vyD1nA85qhRAdoqgbfr
sOZa2KU0AdXdmn2rrAOJCxqgw5f7CBVsnZDcdiaYJXCBiLxEq18w1ktjZy05DfZFORTfRtpIsc4w
x8oVwLnzIfANeHDTADgAQ/bcaTR3p2WlrsohSb2sKy7y4pnQo9vwXBp0LUQJfhyu1HsghXTIlBxb
s6lRvOgE21U3uJrVA1JeWRrYc2p6AaM4FwrEeAB3qcRbfaE0/ztD5C4baIw2TIrPoLwvU+/MAKX1
3G1ICAC14ZyagmqznxHE+v9Up8cpEXCMRm/rR9Hu9Ruq/w7y1l7LmlRXpRvFul6cHR4i/0v4u3YC
xxTNJK8I8BMHetL6PLxnWfjbz56zAc2O77EhjROrVxQFRqVC3YUDl921G61dF9CTrt9wjUKo3ERm
aIrmBRSsBShDoJd2DVl5WgCLhM3GND32EjunBV1xRpJrZJ/AZRVq4MjQsEkdGi2jfaVZlFw6xpaF
H2t+KM3fFnJCXdX2lUDmFiqUct15BMxC3frInFrxQnWf8/NhgFQpBDPZ6iY9A2MUc5isppxuIvzW
8Y4Hw1O9LedRFRpA4U6CWz0HRiBIe1ZWF9XuTaY1m2CI+Ww0WVETH0QIfQJ32wxIFY72hIOLkS3s
1TuOA9QnplY11+dtVPJqxW/BgEIXgecM7mjRLkZUlFzUYrMVH8PoPYPor9GNFT1O5b+WD8aEIo8Q
JP18s2PPJsVK1jnNnfm9jJlimg1P7O+4iak4mjz4P/957hmMNju998+4s/Olf/bZa49Z4AwRw/c5
jH2Pvlrk2HYLJVVuZLfu01SW2vWRZ7uon1Op5VOYnwiNVf9wfJuSjX9m52/78qyGtlGk8RTH93ik
J121Kptm6U2Z5WauRu8eJa1hA4OMGQAcEHQ4wF2LfD8WSO9HTbP8eQ5zaFrr9P6l16OzsmH1/owT
0FHLkW2O2xQIy4uBQY48vn8FpZIZwCzu0RdTsYNY6Oxirfuvcd2UqqnG3U4KBPghncFEw7Zd4m1M
VsQtuKzGcd2BpshJAUmXKCK2AczxGYDJIH4UC0ipYGNic1tT207/AB3mw8ODO6felKO8z+knt6jw
RkTzI92EOYWjxWjdMGaCAotjC1GCIdktcCI3UIngNCPQ49y+JtlbsS26cR8VmKQbY4Y1ug8iw+hg
0oILKiuqehBuypaMgsIlYOIVM4/SGB9SdoJ9SAQUxxvFq2iRqVKqflDFhvsr0q9iq9T+awSKKGCD
Tm7k3c6QQNmL3SIyRe6acmmyaIyLaD+lxCBY8GAjD2WIL9QCWAgS0AgnODXa/HTcoH84LWWrqwRQ
8SUIUtsqnKChECvQuGWnU4n/LA8CiCPcK570zORcdWAOkYh1iG4up9u4iKEx2xikzi14xyOovnS4
//vEQKZWc3cETdjFOEINj/wGbm/7+RCw8+qm9lhQRB3LTL+JJWMnud95XaJ22Mr8WaDFeXnCLuLO
/tqh+xwgzGRb5ALfXMQZfSN9GNhhXusvVvrLSsGSyTe4Mh0SmvnzrqGiMn8hLxt0i5mG3yniSax6
s3C+TvfnpYn6OuVjHXq1FbVxt2HvPXPzJ2Q+EZM6Z44KwneLzJOHIdR55SpW56bZelTUuI4wqgz7
Zcra8K6VXmE3mX4DusM94HzNUA1A9wONv/Je3hyXZrfQLBWGWWvtJCj4TQ96Jq3onYV2YynBz3qu
cUqVv/kblnDcP64jMf4Z9c+WR6DyZRHqztexySCy4LycV/QW+rGnNyUmc+YPW06te+N9fiWCXqva
hFrnn1xkgHpc5xmXCLYRkNFOA6/bb7qHRufGbhYEd+Ho9ukEzms0tKeWwVpcKyNtxobyNRVmBCYg
wmxAl98rI0+QYa33YI56X30Um//z5KIxubiSp7xjCQncTRC458gRFHoWTc6dxMA5LjDLTNtRmUsM
KTR4KoGz8OIqMgWkB2Sb/xhvovaLaHp9ZuXiK7wxqQHmO3wd+u801qH8zWirescwhUzGCrmg2PjR
nWFxNYcTDJuibiVpGdSGJkoBTu3g/bP/fqqy7Hr3b5TqDbA7Q+FpCwi7rS/9TdQiw7Q0jhV9ldSi
vsDabUD8MGJ4YzWTNhXnTZyeiozqAPBUlF/Ccr+m3WM0exff6AioS8FblQ/BXpsJCBZ6JgGmSrbT
s/OmFd2WRPSjUwnEvFNaTCM0f6HFhUOxFqmFxDqRXwJKLI48fDZ54iJC3yT4ybTPOYYX+SoCKxTH
fMGCf9hBBtnf4RFFgt6NubWN88H+1ziCV51ASig1HR+XpkpifruxcbqkTua6wucztbyKfCxJ+FV+
ozhGT0SuvD0wd1TTxIiKybOJs+71NjoC5jtk9KyD8rymS2dVIT3kYRzLRvhshNkKFcqapYN3WQZ/
RW2DYKqWjoHzJrVLlPYRF2ERDbS7WxLAo+RYZHrUcRUenfIwXta1iNQrmX87wG9BwuuHOacFUfqv
l9KxB78IFSl08RJu+3/+ZnJM7m4A3OBgdNwIuyE0hpjwFs8HJ8nSv4WOjAiGHJtNnb0xzVLvWEVE
0bd0raFku1gmhYAV6MEpKQ2pgd6mJWWR9qpub1xJotrM14bqVqrnkBR+whyLi2+i1JXRnmRx6VVb
1RUBGZGBoBoR9ySFlr2JPT5mV9Cb8EJdvRuV4Va5pWMcfbiLxnv76JiRTnLdZ/SVoY0sAfVqd0F6
0QXRxrMjUmx6KtziOEMSOnbBudJQtGfFA7vI6wNCB6z4WURgk9DegO/+1a7xMLNkizhX3STCUP1p
Q3SjCjvXZoaFMaFYlqNx86CUfQkS7Jlec0meo1UOyKQfKFa3RhkLadY66YtEOl+fjjKxnnVlfXPI
3bqcrM5DlPprcy4wc+AvxuRj60GOxZsfq9cTn74guQb2ZQKs46eLPPgqkwzD9w9MY2DyDZdysobX
iQX7ZBhhuggt7y/O0z7OIAe6ScJDo5fb3qTsrQrDpCsWNqn3x1RCkhGanl3dNUqQnmMzvU+SnRiq
VPHl9JWdA7U5v9vEcWogjqhcnbButK7ODeQsMDPypRKKWzNx11DnP5jVlDcqKj6IyrZz35PpmcK7
2Xsvz0DuxF3NUZTUjRhKlx4pbFoIwNOqDSFAos0siKx1pVf7tmCW42v+WMDg4S1a70f/BJ8l7MFB
sntbs8N0uPypyw96LPe6649FpDN00YLYUHrpB0Y3HIBFeRjeRudNEO08VpTlrLDtmbEeUO5B5R7t
E5H7N1Bofs18nS1ScyZJD13bPanp+iECol/bonpvO0UZA4svolRXhoh2y2QeOX7gaJdlS36VeanA
OQzfhcy5ThslPXppbCkkzkLsoC0BKZ0ui4fADKMuH8WjM/R9PyeHXPoTSmQ+zT36bk1x5nVZ2isR
OS0z8R5P7kRXjIWutOMgqynrTT5rDagCdeMSTBnKZ03KpmhKSYWFxih0+wGfEC/+6pFEzzdoEL7a
A136HeVxnr/SfFoTtIbijSMxuc0oL7a3DVPUDeWv066HaYA3Ne4t/tBbMlVxECJwl5HoDQJNDLdo
bHFuXevnw6aJZ6zmVt3FaPfgpTKzTOvqz3leV9itRPKvyk7JKuCJtUQkSqD/pKATsSz3oiilvej0
4ps50GxCEMRkWG9hof77nYlwaoG/1/NajeL0RXwDmjBvs+D9VLcv8vwW7eOS8cfWgTpbQFctUfEc
VvQorTpAhcjhjpiM5Nv2gXcR1TluFhLN8wkPXflkQqxsk84r8g+QqW4J0bps/FMl5ybZp7gLMD9y
cxhQEN0zX8vp7jQROGz0zc4f48681cbLlqNniH/BlExqsmf3ariR5uzOS6unS2EgQ6eHGz7Tsm4y
RvNdGMCv8gF4wR2NmZCGsI3IqOKHgaDoNeodJJXmWJdLr2FoK5Txlq0GOKrOtu9y24YsTYd1t6p1
5Nwoc08Q9T+6LLrflinjbdxD2LwmsH8lcgqZ/SGVOQ/zyyaKmglayj40xGmkPax/N3V8rDzH2Yp7
8sr1YtlvJh2VP7ECc+a/GH5ntFbnXxVF5nbpUZdsx/6JmyOEUA0rDmSbQETlA8ttU3QRUzpKps4/
6rk/ZsE616AXHtTjs4G2jaHOigtrWSeyr0g68Ca3Qm3e5dqkXc4z/shgCQZZYk+vLALybf8nVPt8
gfgvW2L400jTMSdwG0H2e62J+Rrb88hGXogmowGf5p9lKu2E7OoezmSKhDKJo1Br0IbkOs00hjiy
QdCdHI2bc88EU6nNRjGqNk9hXQuZySrcB0H/HJDOYk6QH23nYp5OiS9YpoHKQ+AvzLu8vYheAPdv
ONw3q8F/6UtQWawQKRe0GT6FxCE98MjhQ3xJbR+EtN4s6EFOq9g9LDoII/MUVV1GM4J34qy5Vvq1
ac6HP68Xpe/NVRAjM2gmBGFwuj0J3AZ/y2tuepCt4RD7ysbGCk+zuN5tcWRmvHVYG47AhuntytDp
BhJqwvjc1tNxlkAEbmzrmZtlpI9m9SXgm5QAF7RL3+CBuBB9l74bqSt11heKqQ8OYC+Hpg/iuocC
WU0I6kFRJkKcqnV2py1qljfLU1mEA6u4qaFhnYB9f5dT+N2E/VzyD98q7g39lMKogs9nYzM0GkE4
x/Kat6PmV27nzpZt+RYdHerQT/fPoKApyBhtaHjtPyl8xz8MYLJSASPbc7EnYKMA3IPpZHNOj6Dm
qHkaDinhbsMzdnoCI/YD0/0W7bqd3jBxuxPrAqJzwkX/qMq+JSOwjdmObQ4eN8+k+4z/OxwyR3MZ
Wrjwy6M7DLjDFC92aqyzTa1eNKKGrqAe5nnKamBuqIbSBgB7VpzDR/xS6a6iUVKKm8z/D9giTy+F
DkCz3Ar+MRia6/k/tpesgMFvnE+UqRDhifXr7OwhRBdXQP1IOVHcWOX7Oms/80xigmHBFR/inESV
WzW+XTTvq0iCCkKHUe0OE2vEjKZv6IXEoOc9sSu2P77fnTakFzXpXiERTznMUw3ruIvtUpA6LNEb
CSN8iribPUEJNOq1R/nAK+Xiff0QtIDl+E5/Iv3cX27UakfM+kgadrlI5C6xaezAhMgeSK/pAi8S
uazDSsJcJOakUcjg46AMpcdBJoC+vhPWi7Y3y1Wiv/K5h7y76DfRwfx2GcA8nQOQ+GDOabkYtyKq
Knuymr2hlDJNGFVQrCdwc6jRjTqHhNtGvfqw7lBow36LbOh00XMTcUotBJbN6s/nOL0Ptp1zKkJ4
1GMOvOf/8iM9GltZ9Fy4fn9BTVdMeFFDcNivUPfwjjbl6EcXNxWxwu3NT0vbcYgYN+LfW5Bgg6DS
Kz7mDDCWL43EAvKJbniamEkzcvOSLU+AZ9u2TAydGMvZeedTVcseAb2pcUrRjr5pIoIUI8+Vl2wE
PXyH385XlfH9kuAGNHvBFAR+iCYvKQtzFaCo9MWCzrjZ5oZOGB4iPzCQ29RDjQM/YmbgxdAMsM4f
cy7TZQDNGzVHE3dnfVXD0N8R8NeOSgttr0sdUH7rx1NMSTuapigP000tz9ClF5GJ9QSZWlO4TIGx
CrPn3W+AtmSU0/6lIEoee/9c7yYeuQ2o2FdIhKmCGxgG2rsL4AqS9cQMwLYGxXmJt6RalS0teEVP
e8ZnQDgj1XDTWClERPZ0ZRol6FvZyfrmFrzCZLh6g0BXXPCoOwA3GIkrkpsHlP8p6kZkVvPne/+8
x6HhOZQ5Wuqh9AwTMzDTUhQRPYMgbMvC33/wf0YHFBW6ArtbTItWSk1oX7SXYOCS48yqXUgMHBjv
wfUrJCTIaRGO0deYOSCFGLYwjeWG3fKLXA/QVKSy6DrBjS5IUDtvcR59TGCww4q2M3PgHynn+myL
x8rirEeNU/lQ3ywN0r9lF85QHfNNBUL1rTjXdgwjkTH5TBQ4rIJL7gDddNHS05yO9NTvvAeq8l7w
Sd2dxpeTnR8tuSq6of6bY0CqqKPoW+8y2O6LrPxWy9hHGsKY837wyfS8ysVi2d78M3Z1hfjmUkHM
TG4TX3pp60fbKfmJUyTjVY/ltbcUV4xTxW6pTddwnZLpEZc9zOo261Qb5PiRemol8mAdQmXW78Qi
n2yqWlSQBnP2qeYyU1l8fKsXycKUFLFDnjNbVhGlV1KcRHJTRS/51ywzRX0wVZ/Os9+/GsYhAit5
IW8bVevvyu8rz1xHPm4rnapmBNjiIIcJmnfA71G7moWTOl5ME+/AzA5zibUWfDRRuDgVVJ0347fM
nQyeBhc6j6yfKZ3E86R0kCiTC6TQU7EJNss7ks+HQJLj0l0pelVp8BHIjuD1Q0HOs+53pq8TP/eT
S/P8az8vdhnqxGn2pGukBNLBu3lsO9oyMit5lkcqxA/2e34I5WWCVwHny4wePhYLnfWVmlJqocDv
rdZ76j7bdsIfCpwTX2EkQ1/kxl1hSB70a41MjCMknN679patFxqI2xi/lJzX2pIYDDad+FPMlvEX
hAgfANgIBDz/hYngTnr78GBn0z+vPeBtlfEREYc3lznb6lAbgwFPc4YGYgKLaw8tVhfvfBKSv0y+
0Bnm75WmPJZ1OqYZDpul2RJxMAp9rfumWgmK6yYHP4TcegeD8MZa7RwRSe+s4MIxvA9SKOXBrfdk
rJJgJ7dGz/p/X0T6kC9sZgwnf5VYEExFjl0H25vO8e0Cm9lQHzi6oVOUMZlGcnt0Bv5gZLLtX4oA
AiorW/Hxduoo7dRUka/u6s8dsbdIhJy1CoC211oRFhucS/TAxgPK+SM3lHeeHJuuXNyprEeePHQx
xhvIWxBXZtglYUVseHfggSC8dcjlgQ3GUU0e0E2tHjrPY2nKL/VhANv0RW47J4oSyjgQn3EXuvTh
wJmRe3O4XWGQNOOiNZW4CnkfmU/u5IAB7aesUZT4lscmndskNaORWWXrR1SeIlyOr4uB71NUWAMc
kayggPOx5mL8hjXycpY7piwArS4hgg3g6a3rFxK6nqqjFcRHVwAIKM6YUGjP98tdlhJXyGUaKkRI
x8vK87mqXwKh2N3DVfRVfrV0xB6EBuVGu/fEIHjPXhQ5+Bp8aiQ6NGQ8p3dg/qI+Vp3VQdv3Yh4M
wLLVNwRgYJPnL+HCNoNWZzEKKKU4GVIIIn0HCVB7imnm2o0FsMzVoy3ZCiYGoWwK8ojZhNFp1s9U
J9CGxpcNXlvcb5XlHyVZr+lgOaAxPlCAxfkBzzSNBj+6Ap4qbD4HzWPacXymYx8tHN+iKc/Euesf
cGtnEC7kictMqnj0g4+ByeK+PBbrPN48wQsXq6BH0+pZRjD0bPns8VMNauuDoyf/xPFXzkpfGVfm
NTsX5TF+uM5KCMDNJrpP7A45o1TkEvULz0/MWd2EebMqUAQoHOYeX+WcLQ1sJmaBQ1gio9RIij7j
8nsBpHIQYtiOZDYKHl0U3t0kEipJo0YjnW2gnI5mWbUUfUMqZwqHFdEs64WqQgi8ou/P2fFyfcyA
7/IyF8a2js2/3ZMOMMbGcYyBWlbnV5xAJuZHJMlQ36eYjM15MB2u9ipxV2qbj2KKKkB3h3nMZ7VK
F9GNo/kXw1XB88FGRaaKhxUAjjdLqMRY1TmX4k7PxcQJV0nvF6xtSHQR/9x7xaTN1pCAjUzntomN
xpwkEYxkElFRMSgh8eWpSV+NsBAIXjHxUzKIwqLMRSJ+REzaEV89mSq5GY4VaTCSnkb6IU6Hh7Xd
2xURJ9FCt5LcC5kWcrws4v34akGCt76l0jB1JAMRcF+sJjTH7oDG1ud0YrrVCBVsn2pwgU7D1BRq
IVA8h11Ao09GHfHpjuhB1s1A9irji4djJleMHLqy9u2pzLUSCLwWxOFgAzWoAwOjPpqqOCEOSVb2
JgZm/I4su0f442WvOf6J4Aa9sEHsrXneyvqWjPwf4sH6VvVDDF7PT+4mSGHsc0mdNTVMYlDD3xmO
J8/z3FfZXy/Lf8LY841/ViQ7Ngn4IWpFwXmnWgrVlZfikCu3GxmaJjaX4yQgvuVxiKm+xUhpXSF0
LTVtZG1WV1yXdMrIEv7ReWK+Q1IyKZQxb3vZo6vE0Ms/gB/pqUN6hwKLd1PckAWzfkJYwVY5KfFF
OuyigZUiBPXTEsb63AsTX/2fS1KYqwEN04pJMqYYopwW2CTtgn1urdZcmOHyT8TK7sqQv7MxN0n8
nRLbEcEuMKJLSs2NZwpvZ0F6mCKvFd3h+iF73SDdt+/yWG2rVbueNHwfBjYbKIliwSw4qR4dOsg9
3SuuJ0VONvVX3iUuEfmPwEpxc7Xw029OHH5XQ7WVNtxyy/tBDhnViC2GNgZyDy7uWgVEDG8DYa8J
dAUqKRu0hhBj6wDg0ffrV3u50/jpZ9raM29xFd/5JjOqWLmVVSMTuy5YgImSiX3xOEly4g1mdQdE
mfsuiVGwvHniZ2lLFhmzx3AIhJCYrwB9yiSHUkj0lwbhBHjo9kRfXGS3n1eHFLmP/190gcjiEhhL
fSayKwKR4mPeGRZ2UabiQDpUSQT0gIQGxx67pbP/EJhVZE2Zt1E9H78xulPSTYyVoKNd2ZU3WRub
PeIlUjniNEGHKI3M7BmUY/ZyZLvdtExdT61FmQ8H7Jz74wXo/OP9nkcg77ApjugMdjhFE8KHKvKJ
cdR4P6duVWnYy91c9v026/WufVWvQViMMqq8ahidxZQV22gF8YmKYFAwJo8Y12f2nSQy8jRXmpLs
AZlcxTcDEHpr6HfBQb8fd2Ud208m08t4B/Zt0VYFh/eA/L1Yb59OpSdEWHtbbETpbiUYRgo/s41C
ddWrGmyIDKkXVHyXTcHO73qws7MRcYEoQHVM1ppTqyXViHJWfsopdW6W7vyHgf2FDywLZGCcqyoO
BMtp5ZRFRnBZieuwL8PSajkG7gq7OUa6FOyPZ0ZtY7hTKPezwjCfr6ce+sqtrzoMfq/QaJdQQdcb
xcPb+/r+Tzk89PH623ZScXAxCVXBCG7RHTAvXpEx7ZPBqWlLn5NE8JJS0DI3ISNrjqhnveJFNsUz
lmnZaRcdQ8E+nKjNYQNreHNLr0XWtqTXw2hpY2WTS4ZTJl5Lz3IASDYD18OYl6bFyz++MgzshEYS
wE6uR5z5P5F8+GCITDI2z6bUxUM8SAbXlQYePCkXOF3d1/k5DavtUqb4yBjAw/kYFPbuRHHabGdD
iw724/E5x+OwYFifshh7NnVo7g6kCx9b25NvUKn684qD0LCNfHy5rAzytX+fbO/UBP6JrrBxAcik
L72pVSqvOqqAbAl9f4yQtJyVwPVqa+Uq7bVPH94ceQaah5VCPj/QrNy1mnJnP4dRo/w6T03ERHh5
i2kY3ni39dLDPPCJFSU9XxwCkZbmfWZMcb47c7t+qRzH9C6TxhgWmb4bGye3UboeVS/TQ8ANnn6J
xMiWQEJ4xdnPIxFF3z/T2qUZIJ7wW93r9/T6txAVXiSfufgb6tk+5HBks0Qw5SvWdXCiP74D31tB
FxZKOcoVoTEdM78WJ7FmvFGMn2MPLjARgKIU+SQI3XDC4CDKt21oJr/jzkFBSNA+Kzrve5GIJbAm
9UMb+PljoEVYNazqmxt+uZ4SwdjTbL1DCCbTq9h6fJTObcnmLGAReu2Xouy1ZamLhjcgtBxOm3yX
Qq/CLTPXfbBB8ZdQhECURw+0JfN2G8Qvz6vxHFvq64S7K/YpQTwJL34OtfgMawkeB732y6eDpD5d
l7NQEPt8+DlNxQvIcS4C1lyl+jaP4XE0OksvTu5w7/BCadiDpaR/by1mIRSwCKTlUwGIdTg8186J
AoYceYxND+z+COwyGpoithaWinQQFymPrtw4nZEIjjJOhtiGe0xd5EKkUCa0E9zvIoQYqZ8dT4vy
hrRDtHcXRlKf/o1tv32a8eBx7sTlTvrm4XeldJMOODW/pFYfIKEyQL9eq2sTtiFm3ZkSY3GeKOwc
IXEW5IEYEA4qpekuUQtC0YVnykTlqGmXNR3GhAEE4EozTgzNUUW3Ds1gnVfS5W8DWzTNKYPL03Xm
KXacqSNnLBaQNad5ZwU8mvUyyYRO3xPYGPuzT0DFNnBKeVoTO9MJrT8biEe5WkvLG5ILLPHEp/QZ
bkWsUx5Je48qVhe/Z8XDCPi2M8mQtGn4bbft2IrTJNiU9DMldgAPs85Lu/KPzSzSa2u94Hwz0D3b
HfyyWicq3nqhmnFcaLvG7udBtyQ7NWdcaMi/7VWRQBL+UoCyMZpc8mmgspyMHlLBjIpZcngqv163
hvVsnEPf1x/vw50jUcIy8dyZByrEMzTtvwyBbspRg+n89oF1DVeqYg2968VbgAX+azHuPlwzPJSc
Y2l/wPg0+c5YA+Abxk7nvhbjZL7L8RAbhHogkGvv/HfsvH2Mx6a0U11WT9kA2rtfzBoc+eZJhXuD
JgDfchCISSPTj2fCQVpSIJ697zQs4QM56iX+8bb/hC+FYh0dqhfJxwXDXvFbVwgBgqP4F8Z8j3Hw
c3rrYxcL//e24aiipW7E/ir7Jy2tZmkM0eCxH2EL66D2QV9HQJfRSR4zGKozFBae5abVP1Exf0C4
QnScVQbbAE+Ct4ICJS3uO4lnlRRneb/Hc9jDURyf5pNEyzO62oD1jjEsknGROnMjd38nQIZO8TxX
CyN619Sjq2waVXSv7nw0epiF5zBodSZywuQ2u9eDh4P6cfnwBc1rEwtrxNL4oaallVR5mXIv9AAd
sHlflgQJ3bzFuGD8Ae91AI8LkiNWKQiHBw3N4wcdofsitCONyAEToDgHtIJeaXgy1kCSKDr9HWOA
m3OOmM3WEPpK5O2WTksx1W6D06vRjYPhArmnOw/PV8Uu3yM0vYobfzGtahqjR3EIBffKL5mAPpJk
+Q3s5aOyeEoq8y/F4N5LsG4jfy64A39Q/UsFZKCYyOOZS1Yr1SdUbfKia+CbA4D2+vnE1S4iwEdr
T9kdqH8gKaV0o3ZOa/vMvEkzdp3PERn0N/TsOcrAzA3fK75/mbisyaBboZSGLiC5/fQC6kQ701Nz
TIQL7JgYpssMfQiFKJ6bh2Tw2RUgTXL+dkmVu+oeQI/U+TbzxfrqmlFkloI7bml2gXitm0s+LIIH
vX3m4iwzLr5OQXLxGEFJceRbxJiOv4tn98SHUtCB/GEMoKbYDdMvhKif95+NVRJ4PReS64Arq3ye
gFXq4PyRd3ZxYGaWpmANn0j6ZKdW09bouWEqWfBt538Tducb0MXinoR6e9qYIO/4ThVGETLAdhOb
K1nC2wVKqKMaAYOMs7x0B7gX9O7FQp3zrxiemhURpl8i/ML6DR/emZsvNUqFEEn8MrZ+lNIlULWS
gNbksQqzKE/fd2wjDDErYj0DZdT6EmSRTQkscG97DT2D2PtWgNqjnSM3d9Q1NVPmBYpmJaf/qjOB
KN1z6TxZZFH+2Qp40ATx8qoO65ncJWNj/fHeZWZm85gYNFkphQxQj213SiPpcKcxTh/RSdVAkbvI
4g722z0Z4Dqh0zet3jjvAMQgXLMceQAHQagMW0Kviea5GKODWrIFZmsxTghM1NqDlq80fFAi59KP
Zu5b6K1/uszrlxK1ekE11hjZ7DOlv21CRSiolJKF35TDWz+e9db7I3xuo3rvF2zq+TErVno6LHXD
yVTK0A/oweSST+dDCd089ueBSd45TmwPThmwptPqE6ZxVYDGhTeZAmPow2RY+YFdmByB9D7ZD89G
wxbgWmR49GMeA1GZM2/ks1+e+1tr0QiXQyzny1Zff7dW66tvqesD/OLxu64FWO+4fkR5GXiIFLYE
+i7tYo8EigLpLrViTRn/Cs5ufu2yEDnhqeowodge7lJhnkwZD43flbrseqku+bxxAjXkf/y7mq24
0tkt14/rU00imlFLM/I9hgnU9Aumo+yhFGukXGr2fEGqnOHWpN1dEiTIEhHSkP62hp/Q9MUeRwfx
9hhR8yQxhKjaHjA2Okeemlu6fPmTNHgDu7Ue0BChuLpk1d/V32K5FA87TWF7Js04sj7AW6h7sDG1
QZLTqmqttBH2XFEup5dB/u+iQ66+yVQa9M/8FMlA0sKP/0bDrkqyT1NNWgK+CyaPEUCT3HW0zKG6
wuSaT4tmrzaIvJJhSM6F/cBEGalVUdzNKQfYxVJV/GhhrSVtp5r4n7gR7yqKsKsBQFx46cJXt64C
YLchIttP06xuAp5Pktd8pqm7f3YoXiAbikULgem70yfCmpeLwBBZcddzWbHoQ796dreuQ/Mrjr0G
z03wtTHmHIPY9XtxgOyODcaTvpNs4oKM5cpfukarXJMEoYg0zCWf97mCeHWQM6iioL/zILbV1Jw1
HK3XrqFpiXVyDSfCOSv3pmOPHL6XIH2qTe0Q4HDi5IY8b7Cb1WLZ2wnEPnKUBp+X4tVpRWFc6kTh
gnu3ImRqtSD1HoCEkFW9MLPblYEk/ad2z3cQDYWbEcds8iVpeKMV57oXgkhUtrys5yaHsQhkE5cW
WA5P+8Y7ZV6F/UaFJmpB6WsT75ONFPeMGz3o/HrpEmeM5pjyghRjYFgf9Y/cUR3GdiuDp/RKHaJV
3i2rwphfv1Swf7ZqAdmIj4zdycMl9Nv4eWVpjFLSejQvLY5zqRS0QCsB6bcZrHn5sKEgxuEp2vTQ
KD6Vux8OPmA0tvuQfEUiSC191pyc0kzPbcdugvcxQUl9TqYj6MVWoUwFNBEVSI6M+tBVG27rUQvN
94QaknsZJV6lDwKIph5J0ZteoZ+E1gVHAumZSr4neVoyd1qrCdIMjsFD8LlxQ1Y/WjFMiUppj8td
T23SxXQHHbhoPKs0W+Mdq/gXhMy7lL6v4Z6t3wMyav/D5pUojpUcrsH68x8SDTo6HxAHDqqP0Kin
Sx5stfWlHGWmtQJMZ6UaBMhp1pJMVltIst+U5Ll/L0q4N+7n4GFKITaCIAWt28guMKT0X49mV7l/
iUgcN5uwWifFPYl0FgRThchOtxN3RnZy8cVhFbT4quD9JmqamAOVLqeqDHs66VRuWmn65nPEYqIP
AGqCtzk4HkS9dfQI/SMbaPoUqyCjJ/thmbiIK9VEKjZ1j3Rqgs++M2NGSZbFTFjDepanRJ7YL36s
pRfpBG2/bVAj7A1bVPB5dvO88SqU3Ap+EALGsaELnw0/WH2vUSBGegbgtodpTlhDJjogWO204PUP
C1qrn3YN5b6PE0PaptOpSKEpUbJanlvTa52a0doAxIGCXcyhMZr2BsJRpRa87zBL1vqn79RRQ7Ib
K7eGZUFwtxGxwizpScL4cLZYXEh0fcElECReQl2RXE67MwZ2DRa+/AJWQltoidEGClAzm4t2f65u
gatS07oirQTc4AkQ+PmGlAfFTGT3a9q57aIiUMzq0CG0dUR2asxN1OPL8grC01iKXmHZyvw8lz/M
aJDKKFk2gSz9RBqfh+WZ7KvbV7xPXt1ZfMa8FMwucAp3MZ/qO6l4eq6Ulz1KBE5vlGaBYbLABcQ8
A6dgg62ZaRFdv5O9SkY2BTFyCMEy7w7K+1+oNrCn4QM/VmVbGgn8RwFGlz3B7VZ+CFGi5ovQghfh
+IE58lXbMtJMzFdr3YHjV/HJsrbc+fmajJ3/aFdcYj4teKVmJp6m+d/a9cAg4YeNvbnx1QnV3EQ+
RHTj8uMGuRbbuN81Ze//nZdOx8YnO8hr8NDGKjjm94em8kpc5ddrByz1PtFMy48GVAqBiDDZZN/V
20dUsBFtbypFGV2AdaFJfIi76dfpXrH3NFv0K1x77J116iqo82DgCheU/xAU3LQWZNpvHHQEXlFJ
NbfalHk0FLCHgzgKKjoMtsDM2+qWKjD13d/Xl1rUgnJ+5EGiMEzsU7yinj7RHICztFN4RubQYYZ3
WryE1XkxxZQvCCsA3h2uDILqTyg0mHwr6/LVA4FAOEMLHLLPGawxhGKx1vOtbf0aIT16eqKD3qEf
iESwV0P1UEgcK0eTvQiM7tJNrc369kaQRwI1N/84HCnf8U8i93aVHRxm+ZXV7z0az4Ik4e3CdZcR
jcN9wgPpDs1yuu0EaRqz842fVVww5ranoEMdORVjooWHeqgVzXzLlYHLb4vsUFurkollKo7qpzIY
Yk+S7OeGP+prZFwkikr1oZNCNHNxRL2bEp8CKW+X+Esl3XR0H7lDzT+W6jvqzG6WScLHNdrTP5gi
SjLasR9zSFJpm3C7nxx/0EZKFSTE/jTwSmhmsOFXe69uvSmmcm58ozWUYfLscibEPkO8fEuIu497
Y/nnn0IS5tAyWlqQ/Pv/2eFA0BhNGoCnscYdCbBDetEU5VnXd/Ykj1PmuD9TDy9s4iUHqtnxM1Uy
T2HyglcKcHLBQg3mtChqYrtnrMo0O68w+OiNzJBa7FJKRbAxLH5iGf/2ibDCQuGDCT6HKjvXrXBD
KpNzIVskar6kFF/lePeNR+TyCG21596WRyDK6XGJps5XxM0SXdu6y6Jre1NbV1y6vSDTmSTnoaxE
o4nSREJOxQZfrBTg3dGoDfOeuMd5ERAQEiY3fvNah0Va6MyIfo9ZrpD4eNVcVNNJXEGMNm2iwyUt
HBJqdslrY8oRh7Q5Q9EPiVMtVx8nMCewTdsLf6H3Jj62lGZQJWHYRos17RBWWB8Esbl4HtPHhnnK
jbaFZQWmYyUEFmHdY9OklYjUXT+6tv+IEkDWnUxsCahbjyGIr+9CHcfO08zkxxnR0PWVPrv7VPID
ootinbz0rA9c7+lGa9udTBPqQ3iTBG6rOs6MdSsKzsMvqMPT8fKd5Zb0Aoaif64Akekd3LjuYB58
AA9MEcXt91nluHABPgesHF9JZrEVvIJOa/lRWF4QfZdCDT3YLcxodDu33A5dk75/V3D/6jL7o8AL
kfTsRIU6SZs5H9ytS8eevszzw/DJgCWjgO5khCP/Bcx1x3rwqa0H7duNCm1VYr0c4H9BDBmzPUgU
4cIGhJqU1ZVI0HcHkS0tVlCfdhiU28lUg7ZPsEzfbxj982LfDIYmXuFSNvbzUegvpsx14ejjhJS9
YgGAz7O1EAnFtfwdYaJxp3/S4W0hImfjjR2Ibne5IeIa7uJESh8kaOZu1ikcyf8LSw3qyAIe+J5O
XzgUpbAfyNPT4RmSbPApnKJ8jJAf4oO7xLPwEvYKf6ap+NDPlSSiY2k6k4somFRadtYA8Hw1UP08
QhcfSCut/FhXolo6cHn5SjBfYlN5LVAgKUyrpOsXfSdzaIi6krdRiyLseovEoexUyKUzd5kQbYJ+
hmAj5B0+Gb61/KcbFnwrGhydVMiIjtzNe0xuqqVEdvK5XIhyIKLbLl0STm2qRbaOpeuhbe92Wy3q
D81Cgxmowz5WLQLylZuhZ006swlVqfnXj1jvL9zrL92zYn3+2DiOC98NUGZW3UHkCwSRPNi9eSst
BS9OEx/mL/XWHzEeewx4tw27b/baJHtFYBCCyWgxRLPBB7xWqA1z8G9pjFZWVvXVsiG9b0cKcGBL
LqI+OsbzOTaJJCPzwYH1GUdAmQHSQyCL4HFiI7HoUf1lMRRrJ+phLV+q5soxTKfMEw6J/aKS0+J2
C5bFEqPN1B6LQMRttqvBurnmzzmcONyZAjV/RMzObH6+kgV3vuhDC3xG8L4bc4TvsIY7DZTwtXCj
0Hxi2Cdj1Kf8UxWnqOW7Ore4jkk9iSPPk9UPJM/woZYRgpamO0LO2aEQwbWY7Je70G91UQ33Fd5J
P/WuTgG/v3sCyREM1SJyQzEKiqG8dWpyDZpXgYg3buLyz7BjXxFSU9hAmojfXHwXQ2Blfi//GObl
YfyVyqkESTXeH094Rxvopo7I7SfmcPcAXUCyAI5b9FmDqCS3UOcHKMDbgVkJ9IpE9cJNKIcnqcku
Fkm3gBXkXDxjhN4F509F8+wMstoQBvN7PtJhl6F6qZsVE3h61d+9ZB7y5NcYyTFJCYiVrU1BiYiF
HglI8JmFkStJLSBrHeAkKZbzqrh5vLvHeIQRMenx0ioZr33l/S4mzYVzY4fUbRx1CMJAZ2SSIdOJ
GuSGF8cKcbZz9Yj5A9Ude6MO+aoEYvaegYYGp0XryIN9j/Dpi7R39HLqGr6aBjgKPU0pE8jOnFUq
Il5klY3Ug2ndIXdzIhHmsAK5z0cOR1CRYQgJuYDnxmGHZpKbUGqG9OqD1tQbli9vQCNAiCj0UY3f
NcMwpNEL2gbGTBFYXPKRhXITJ5dRtb6jmxpHVxexaP6o3IoE2tY1yBHnjGH0n8Ha+5t3QOyz+GOj
1onUqfJV2V6puI3rbYbi0urIHRSVUPid/sFiMUKI1+3vC8RIl+1hVWb72K2+E7KfWghcFtX8A0qF
SGkvljiVg+qX3DQsdQ57NDc9oY2i6BqPOPcvAS2dYLufL4zqpXGWyJcPYgqeG4PNqKbKcYq4YSHh
H5sg8zdqIigoJ4Zxjrh/UTJpH0k+RcZRpEVFoUfKEBWGvktb7pOKgyp68llK8T97GQWeDaEg8uE+
rHBQnEo2uTk88Qg1kUSvIGv0cdcazXMhrVE6OID261gi+sn/KMuo/qHg7gjzWEha8VfY7vHfOnrB
+hgHolxh6a4nzAEcgBWSYVLeT7x8z9oIWxbkt+mREg9YkJoOiNCFDB8oN2ELTtqyDL//J6swnv8F
JC4verbVSZW951+HD67TT5saSFR3RY3xycT0ZyubTpwH8yp7+XcuVSpdQOJX/B0K3W5k0UJozrKA
MWwacz1COn03NZ/GXzv6rnR4snI7dqJQpGz9aFvWrtJQJ51dj+D2FpmQH16LKqexC75saNYoRVPp
5KmRFDvBGsfor7ABzUsgPKDQdWRiCu3GNDkHXAA5LU2NuX/R1J87gb/IaNUeI+ympAcUwHEzNP7o
YAd0OJ4eD9bkgjWRUfHedg4ZmF4ts8eMPE+otftXFiiHfYxp0is7YY2fIPIdSKdbWbGwAoUXxAm7
iDCBUjOYJrCFbkspRi5IHQnL7x6aqD/a4z+BJklCW/HqG2ZqXzyUtKKij9hbMXBqqcEMDJDLAEUW
pUUvy+o/+S9vXw2cS/qjxiKfF/F5aSqNv8+GO6JYiYxkhIq3ZQ23n9gSPYjkfdJn13LbKdRMuwnY
Gg0cwUjk7CtaWF/n5VBTA3cwKtZLT0+hdVj7IU79WZ8RF4IcLI2AuYl3l6SZXgvoIV3NbT3dlaNr
7De7/mMUDryP/a3hgWVjQf7z4nPFRAHt/PLozW9GH+zV9BktFPuu+gw8UdDeLvmff6fDXctVyv05
ZFarZHHZnc5dVjEyW7qlKd5fqZx+CoY6TD4o3fRmlB0nmxMe7WRdV1YsMk/JvKc8SarYREFUlPUB
gQW38U5AMPeRnxP+yt8t1vjRnhWCjysbWPyzHpl0ARlZaUoWR+rXDG7CCn+D0th2nW3ME8V7XoTA
9WP3lcA4/g3CxptI8mvBO1jnGy3UINDdAuGIjdBgAjSZxP3nOrncguiWLoWefVbs5ps3AzfcHYy7
3YF5rR2mSrNf4eAAFfBHIGIEh6Kt4I2lhFno6SwEdBWnpLhpIjWhv+4vRDJ2CRyDHonde3ZRPtZZ
tNrt9JsaibbQwXQ8fxztNOryKBkUS/OHrc6eSVDFRdM4toPpMjjPUAQ+QkF991wTlekPzNjyrgJf
5vs9g13O3GrY8TOcM4rj/aucaHKDHa+wSIJ6TvzehNxENj6ngj3EM9DaMwqy8W6u0mA0X0fUvE7Z
GnNCzFv+waZdrU2EDrRLxVSnkO2Wyygr8/SxWVsAaA58ritxhlxen3rsBzEZXmKzNa/xLJ02IX8E
04sntZ/bU1syrPOLBFkaZ68fzKAlaTGLYZ4p/az50tJvbIKJJ11XQDl/uhAUxxWZrXg1h3UCsw2Z
z8LRKUjNdv4FtILWyjkEJurD32AcdxAal0C6O9WTFEyK7HxVE1Udi8bDssQRr4hoTJwXS2+mONOi
/vmelwz0ZWoXpvJ1z8ZO/BlN9IroX/bVbY5phKpF/KCqXTEU0gtuQO4N5aMsnzWwwWqcveaXCKBq
jt1UUKgsWRbLMpWAPm4sE5ZRE52AC5OJuHZ0pIxXX7XMeJrpIFQmQ4SOAOUoRzTO0B+43fa5qHtZ
5xDTHWP3hLWB+8PJBLm3r6iVz4RcGmppVu8wEUGwm/fpn29v6UttjKMNkW8C3VTi8/CQONBK0iRK
WCG6apqVTaVHAO4UvoXyIrjxUrb/Zj0FnHcVdZbQw3QDJGUxtVWwytBV/lKw3gvp0x1a9SmbmUlI
u5pdHET+qev7YEP3/ky0j6BMUYaMJPHp91mc89/+1K42xn0vMBy8DaFfEV+zar1U8ZWEE+Nmv/t2
AtzSG0gH4wE9r0B5m7f/YCa2SzM7zPYKL0pVuG0LaLA5EP52ONqSDr1lnhBZ9n99ClIXSM/2QAit
XvSazOYdyaTGQ/mBs7zw8PlD8X2j0bGOQJKvrJN+eGIPcKwDU1VLeqeMoPg8h72Uaxko+oCUYbKR
sm1njF1gponNiN+fHXWaP+eFCR9PlcYbjkjiMjm8IDWEYPqvLydzNgP98ZmHkmtWathzv+tR+OhL
+IlcUQ7BovM+JlwDci4CkYBvwQ0F9t/vhwGiMOp/Gt7JR7sN59AIHCVv4TznIWVIVyJJCIApKVPW
j3Blc+B+GDwtDM0EtVONLTICleV/0oF5yT3HIo0jqLB+8E6Ha+HOg0+6CdB2LhPpKv85ekdeiWM+
ddiasOoLSFKFb7vxFmb1G1otD0UY7nWMl/6v1vmHtYdx8YthxOJRmuP+MUS3snIQgFJOnfk8YrMZ
VNLDdariDW+PkR2RYBR+NaPZX0br9IDxA5ssEEBrJEQwQ0KnRVNK418tUyz6dg7EYwET9RfquXxR
0HuE8/lEgPhkzdFG5mCY5FH+5OXPASDdtV3/AZhQhTUHFOLV4GgWNByfXryB/yu4iukHjJ/0uZ+/
T71Z7u0WFSD2dkQcbNNvMNAV7nmNLtrFm93z0mZ2NTsAbuNDHVtSoY/4G7ee3U2ciUF1IYpwAZoQ
sjjJxD8Aojo6JX4A+jrTB6jclHfeXEpBN0K8w8IkNToLDzd8E8WdjApf8sniyHELutHOzgMfSZne
pTLctIkML/BsJZdofLagTPIrwQ7FtXBPvQiM2YglVdSOmG3lDA9CUQBG8XCn2YaoPC/XmBLRVGBf
/myo8+fDm9XW1eqk1C0xDSbljxfiyha1R+oG09euxEVyOR2AHE1s3pEjgBp39j+nIw9ZdFxBhf4/
4g+jkkR3WgC0Oe3q+VTx5GKo5E2ZPz26anDL/BavoClUpo3vcpk0PG/YR7GFig0FN/ebZ4KHlxk2
cCxaYdZr0wpLyR4bKFNR+por33at3mFvWcnTs06WRFyPRPHrTBhLPynk7SWpEkbWmRy2LrLl0Htf
SGbeaLEaYVrVAJ02pzBKkxcutTbK84OwySYvwQAxjem7gI+sJ+Olg59xVFA3iM0Q+s4Yp1mY0dXc
FtflxsusSFcHbjzalLvzxpXGdPROCY2bedmrSP76DZJCB8OSP2ijgsmqeSIbY+L2ZjSu1rRPf2pk
O+E6o+ZHMiOXGeXSj9M3JXBUip7CdZ6THCynHmR0KuSjmh3GvIQwdM06nrwT3POxY8Bwtlsxjac8
rsXGXfQG43Uf39IOs/PUmOhHaQDGg0Xty4Ky/46TjczHYJo3Tequ6HzGujqSsWSc+wfgZHfO/dBs
s+lQ/ZePJSFcRO8DJwHzusTB20alUcqd6iw9ZnzHEAIDyhvLP9kaKshOmcmy6NYgb5f9ZvHLmiIW
+a85Ikh9XWJe1EviSjgG0/7Ojftxjk8Leyh7K9Wn2rSh7b0LecOPDgeki9GYZ3nkSpFKEwM0P1mm
CkiwUQLo6IrK4GEDkAN6k+GZhMjw2lhydOU8QM0hc2e6VfR5krq2Z5Gq7oJ1SEpUKzHQAQmVNnd9
rxg4TzWP9hBq+aXDbb6cvG7GOo93lFTMjrp8cLyUSS8aGoTWRa+b1AYzrrx2tHSOHfQQ+Tx+hBNe
hBzQQHCJQbYGPqWcCprws+A4OmQKr2FfJPpJBrzyhEawAivDA6qk46SPOKYEe43ojl3wWWM0jDp/
+JWz6ylACt2dF5iFegjnw3JyFwwpDuH+YRbzDKLVpJGVGYVgpuUlaTk3dVlgbPSOJU7OgHJu7yd/
yHUbmeGc1Vcq7xwiUgXujf9uVfuVQ0igXj2i3kLy4hxJs3/YQ9yalOwi/qdi+hzNCyo+yf5fMjvn
sOEAHrvsBAGP1dYXhT4unzkYtxo7UtLu+j2mH4T733S02LEnvw2kkN0zd3wSim2oqtIApY1qXEm6
5TVz3ZFMmjK9aV4PBv+OD9ceVQUeEC4bJPa+bWOzW9iDedfO4Fch+lAn04ArosrZpl/1RyqkhW2t
AgghRfBzV+Q4J+2VFrTgSIa8mIfnZ0yxOjxP6IOp6zfRnWZb2znvL6qHMQlkMqGgPSuQfbxCWahd
2Rr1MWyNi4h5M4RBuy4N+OoHuZtOlsdOAgA15ifYo1KhuaRJlKsMBqJ6N2ZD6z0NuTy5k1Ho9aQ5
0y89af4GTuqApcjtkeU3arwOxFzLC8wUiWSp/Y04l7uy3zI47cTRVxDO5UYpzNOyitpCs52wVXoc
5WokPe5sfTE8vJUpp6JkGZA0o16WxX6Q5+b1TbkTAOIROk2uTAxbxkZ2lD0ccVs9016ugvc5isfM
m4kgZB0Akm20FdT5LWRf7ZPXzplmCnhLbshpo8kYxTpz8XQj9wWCGnZOGqQZB57zzSSLcNNN+9wO
I65vGyikiCBJ1qhAb74b1T2lIR+47OCfFesL6CEPTvXndRsR9+5+6ABlcVufcnEPoMUEYhEteYWv
SmTnIlfwExGz405AIkUk8kZ1jGUvZQSB1XvQjh1SjAnl8g+U50nerh55iiyq3mUjZcDCZvfjR7ao
gewfZPa8t2o/2m+QeEV7iJZBCCyHfE71QXflqesjGluFAZvloaCN5ONdzwHk3egqR9LioRpujMsS
YnEWz7lkxy+fHsOetUoriO/DWynZ1eBYQtQrQnPzcmnC8PV1fbuyO344t0mIQoLGnCGu43Eiplyf
trOPTeZXv3t4b4OKOL7TOBI4lsq4AsaHHIg3g62Cz1tIVcVQAE63dlFGD1ymcOEapAq1qJwnvton
FKKbq8zl4TfsExVzotxXWFe9bypTLGmeXuwIHPGBdYVt4tD6xSUTOCrsUJrLMW2r9NQlxzSpkD5U
YIsDfNVko4hhKn4Ox3ztkRMSsdumkIbF3U3sI8wiSSCF13uYdVjcWHde8jimCktgb/Kecr6K89kE
NiHM8xSQ9qaYd2GkqlWTIB8tR66mGMjzRl7aQ0aVr+dYoNzWasL7hgEonfXhdLNsbCtcpxxxH3/z
lvONvztaZulbrcRDdCzSMmHyt3pIxf8BKuD2EfaINyvF2S1yScTToOt4kyiWm6NYqPKo+kHpfyMF
nSjvBArdoxMynqRDAnZi1+H2LctV8Bg+JL8F2fHCpvL8v3qhzRdcuoHqFmjuUObUVK3nHtOg+LLs
BRQhCsq5JVBRL+9VcqyDpoGWshnEXkyT/NxJ9uwx5DVE16VvhA8x0aghrK75ESUbnRl6GfMd1EWc
OQG2vRPcWSfvdcUsIZ2qS1K+LUa2fa3sXls2XSlN7TRZYLs2WkOK5TDzF3UqjFN5i5Nsk9X57mWQ
Y4aWZaQ+PqxjZND47EWifaVlFsInpVHB0KCZVTQZIqgoWfAx5XGbwQ3FQXjqmHL1zDvM2z/BonxN
koMK8qPJZNr6PsPj8auBHi3S8Q5I0yPA0goX1PV9qhyJd/0WcsC2PAlbgrTuG+hUMs1ruBJY90L+
NQiZjnrgsCyvTMAs3PN09zssBVVnfnp5gghGkAqDvXDKA7EB0vzvisPBv9O/WBf38oTZvQ+awAlP
/nc/Df7k4jf1frakHEGYHGI57P5U81NknmTXmdtIoHFfYDfw3ctxZL7JX2ERWSxJSK1uITrJiJHN
fZay8qIqZDKva09WZmlZX7lWREhkyjb8L+kLf0Aos+nvSVpWM85wZ+tTx3LQTYBTnoCfnujBLizW
R6rRMfJ3XmkJ0FoI7WVw7KCaPdyYLZljfN8xA925mHPZqcB0tOJ61h6BlxCm+C7oYiYLkTciYOYR
W2XCXxldm4vZSwpwK9W37JJvv/Pj0xNDrUCWPxviYAEwIND0NgHFVIpC5JKEtEmoZyKa5DZoUPHg
VnuRafc1ZYLUK3OvM2Mkiqy/+lw0tRHDvyPYNg5CYoN0Xxr1KH0uHhfvH6fc4GeaLE3M7APtbPY6
gv+R/fd5Se1kIt85zfc8Fsu94H449+Mr1XBuC9K+BQptzTNIXsIofYxYiOp2Dnsrx3qpznvqYXbz
6vMrZSaXfptkpUlAQvpfYaz7gzJWFmiFMIhGoLwr00lB8ckisaGIJm/as9Irsubf+VVTFZam3eZP
LzufviECj++HeKARI3O8tf8ypVXX2blh9woAME87t6WXNv/gRtFtu+qESo6SJR+IGXqRtM+H3zBG
lHfHKOd19FEudGym9ItDz8iZ0/thBgwlamt0q0dXYSDgWOXqym8RkTM5+hCpKujd4V8TC4g2CaZC
QDbEQQkBUsqmua6V3+M1Ga3XZEAA99AKqT/CTEaH88zJJ3JtOWwZ8eu0cE/J1UCaAMf8FL9TlTY+
lU9ln7azqc4y50IqVpw6vBnvxu1+tS8JUo+uyuELPf7CQMGsi3nwj6bByulagzlFJACkb8Ej429X
TTtUj/PVZUVI3rXQXp9GkS6FOyY9ckRY50R/bAw8jQbGw0Kh39bXXeUztRBqDHTEXV3xsWUbCtJT
nER6b0EJh0CmbneKag7Pj43f/WjugWuHsL2gkAuCMt69nHMGBcVbAFU9TybBBP77bHmOa02IR6AI
aM7h1hVN1kzfh3yGPNlkSqVaX8MAw7OkH2HGE/aB6Lk8MWNFAM86HvDsVgNMmE6etxX2eUIQzMjP
uRZ0HORArZG7TOcorwEvfAek4U1oJCnFEiDjKDezYlrBVt0c7ztMAvGNbUsGeTgKYm+gDvk2aEgr
kjtDY7KK2iSeB7QCxPD5UiyTkuQWukC1zw0bbkn1XjIEuj0bYQxpAi0ujPsgtBIdqMLbIiHdFJCf
Be6IvmFQrBjlScTuFlGdrkQOIWuwldu1XxNYejyucfot+UfFSSpxSNV4qEQgZvEEzP+oIyFYDe/R
wsdeH1bvPlbdGlwj7zwXmWzqfOOLIbYLLJ6YxrbhN6k3ehHyaGjWoFlQZWFMsWMHyJLfO29fkTzJ
lAUN8Ogpd1ywccyDHwpAQyrzzA51iHT0mM9ph7vtpMqtycX0wgkayqIdFbSCay9AizH8X2uwL4wY
qZ00YH75jW2OcUZ+AB3hbqXEarm/PYvB+uktuXz4+Nk29VHcLmuy0/MF2BzqOymyDzYHMe+dPz/r
D91tLaQKiaP67Q/gXULHQ5vxXUleZ6LvcvTGfPsyM2qwg4E3v3zE5+vCdWwVHNU8xfzth2hX4zYu
8Fa/hdKg2TTiy+RfDFMjODIYEe6N2XuCADvdJAnGad57tUBLdjxvWpEWob+I0R3ho/kNvcDikk7T
Ulh5BcYchp4W4CqR3pe9IYv6Xb0DF8gm028GiG1WyG5yTE3ZKIRbzygBRCQH2PtM+YAADPvqdC0s
bh680DxtVOW2yog9fRafPcKr7/J/d0kzBzQarkaob9r4bIVuAg5WzW1//Bix8XrKqXDRMJKjDy3f
kAGFom074TR7HVZsaq+zcNjNTIFN7bBOyBlcwR1dFw7OThqwtjAdZ7EzdDXbLBb3+nEmVX5W+49E
t7lU0m5MR8omlucvEFMOrCL1EpUwEftN7ME+UzogMLaUAIWf115i79jFZPvammMU44yaQmfKVg7z
tiDipE+W2i/LTqJ0REb5QpJnkRTO8AircigTBPzd2qQy/Fbzz3k4L44Jkjl5NXOjGRLg8YDO9v4v
RY+avDRX4Mu2ZtE5beg4Oul21rSdiFjKVMpJMsOlKBKaBrb9TL5Z0jKJiPZj//6d9n/JmQVxDdHD
G2tOclEJPjUIxBeudF1CIdS14SbNKHAkb4hBpOBQTmaUE+n0xmW1+sEAUDMIe68J5N53Fi0DP0xC
OwYhENTCL7q/gqwy171eOQ/v3+eyEp8TIFAG8uO1OW75paQPju8/LkbPh8lXOlMyoziBE4a3mREL
pB7cSfg4FgMsjCcvfITdvUzTCl14JhMns4ce32q9TR5YhzEvd3c7RMt9ToK7LlciErvu35X6v29P
7sIXMTO1e36UmaixmXcxMPRNs9AucZMQRxnf+kij53eW2+5mqkgGGe3wktRDkfNs+plQ9sxMTFqE
CavtkQna5cjwbVUw84Mj28PbqEJnLyyNpXoirnyV2qFazSzqCaHFiK1UheiLgLGImOsqslm0SHS/
WaOrK8SsDOmLdI2koh9lM1mG2bX1FJRTcznFHGQmBRkvLOk38qsnp+W5B05pVxdSgr5kun7+NfS3
PiykDwf59LtGFYNDfCg7Own2A103ZBT7XM08BNQM1YH19WHUDrQRCYrWSrU66iUkLSqVKfOMh4i6
XOcoIv07xI5yOAcUZNiFoGOigegf1uKAsNytawebuMNy/UDvLUkplSUk52VKJ8V62+tUE1NVvPQd
bvhV1DDWOwO8ZgzjiENdKQ9NVQ0Qrvx35MFhMqRe2G6ENX2t2crLg04b2z2khtpvwxPjJJo/oofc
2htKt0V7qCmb1YJOA3zvjWuIi7Kx6vDotyT1baPWCwkX1T4qzOPM/VURPOClHewbHHO8LziBGQFJ
WKvA5Q2dmeKveXVCm6Y0k05Vg+Kv5kxV3OdNKhjwS40lkDk4SYT20mpLlm1M1DCPGR6r5jfnz/Hd
YTlYilWCzRVr+ygQDHLA4w/kupRADPHnjTEbPF4jfsXoE+TFcrhzGybPTH3jRD/E/bJ0/IWeW5CZ
ETJtpCq+9QmUzL9fT6aNoPmzzUg/Ex8U8N+CPSHyBoeiEfOQWW5Yi1rBBK6UOB4yjeR+ECiAqF1G
ojVfCKEs+Qsn6fTWyAKMP6ZH6fkTPEZJOB3ifMcKuZaVk1jccz958bOeupXq5Ods9+6D/N0ld6c2
XSBtypdlEYJRnVIvAAlp0ayYZeczhZ44ImyFWBsdzbrLU0WaunSkNOAMHBk6Wcq17ZN2OoNwwFWw
bwVIDiPBVhdQJ2FggIkj7lN2R9g3H4Km/VipJRS25RcBz+ujq51B8IDlIY1/3tB6qYpZe/qx0gF6
SozeTZyizqnNzAJyoeGj0K7YIgSL/cD3U4CFOI/pkhWrAq0//KxiO4QAs432LT6u/zGrP6mAZb/L
VskEPdQCQzKl8ysiED/NI70ael/qJTyJC9DZOgiT+2aGzC0+VAz2SF21joMLWS7o2UzrTOd//870
JoWzdxEwgbZCyjylUnNjXekeFA36O5PMnrf/qhkKxwdzhNe/+ErPMdxrVvNBpAFFV2UeQM+rbWjb
gXX17zggxtn6ifyRXJfmmQAp5v+SpEomyNIliGoUoU7QOXz1O/hNZGL81r8FJeld3WnoVeHGAR/9
2G4AlOBvlr5x51ai3AStRLWM8yJOaPz6DA8Ya+Ch2IZ67tnu48nplbonXF8XCSejT7zYJrZ+fisi
Ow10+p5SKtYp/VlCYRwvNmvlpAEK9748kAF5fSgu39/C7eaR951AqDPZbenxYGRYpUK+T8hcDP23
AeWYpTrle4ZbvkMSVmUzpj9acSlu4+QvQwUJqG1Nft7JVMQLhLAeVeCIViwGLzss4QjaGk8+bbhx
m/tyajvkV+dnusEIrCYxKtf6kiOQAGgbZCxNEf2nh51wwIKwK4PLIZnG7uoIYW1PN2Wo2a0xq/++
4vdPOS/lWFPjiMF2uvOZ4E1MYHMZWk4TA+DtUk/fTUUqbNZZWQhC3ngxdOysNKV8hPnk50OOSg4+
WFaM3h/e2+SbRb6N4Y4D4eg1VCauatgACJF1BlUXOOU2F0QuZO+U4NtbyNOITDEw/uqp36PA6tSf
0RrqTdMReYXedPpxfyZLo6ayjp0WzkgHNGPgkR3zQThsvoHGSXIPP6xY9a7u+oAtShdZHALdJB4b
Otc9yxqHjRTGMbAmqcTu10lMPgG878pWGq0ZaGr0cMFS1n2JKx5TDEH6YjZRkX/zmpjK2JD5OxO1
sYq8wFaMNwVuLXYfkaAc7wuua/T5yqgSMp4vFP81RYkkrs9n8KzhdNO04/SJosc1v3pToT8T2k4w
FOt3U6GrKlCN2nnSkBS5R/ZVFIADAHvIyWT0pxeuiHO/Y2Z5LQmR8z13MEM3wI+u9j1/ir4PVf46
X0Nd2lXTtxPhG0FE22wARJlW+CnSijGG5+qH7nneur44rbU0SlyHO58i8qpDKlZcF3kX3gi8lDrZ
3CuPG53aqLNoXxfTjkwxY3k+Vvm4E6O3SDa1bgQg1k/ummesSSY98rQ690qp4fey8RklH8ZoBzfG
xBhPWcnOkKOuGAfa3bj4313A8KwUxcuQpBfwsoGxiEnbqQQrJLv9gooJCjZVJWnEKPIzCvFTAbND
d7eqMLN5MyeCdKIgeFHLGDizCa5pNGumxu84vz5th7l0r4Za06xxrhDR0LSgdmRs4UgeaDU+9Rda
L8xgSmmeCDXd8QS40ICHL05bqX/Wp5xg0xaTEyi7avECKCwbnOePmbu7CUH68L0DjFUrV95cn3N0
8ZWA6sMMyZk5Ggbvlgkh0AXi9b+iQiK7h/YZhZjBBWsqsodm+BrSDTH0zgVkRQHXSLmur0kU4Ooj
WcEEXiNo0QlQgVuFldFU3ZdqmqHbw3W61hV2+rhaqhZqyn7pg5V9ROB/4QYdTp2r9lAmjSZve4Fp
FA17Dr+4pePZta9lHVaEjL9kWS5LcdyowH+D7GWO+PB60g4u8OjuPjBCu8tC8A5JlZRyKk01uRlN
BoETYT+sl2GYjgia3QqQM1DA3x9Xs6PjplAPjZ/Fl0AjuCg2BISIdiT53r3gruHCmwZwoxKBnyd+
fK9Y44SzSccLCrojBn/uHxh8PdrHFS8AqWBPBD0+xEjWQseVenPs2hz89NnRdDbVhStEnkSHmy4+
p5JJIE1edUfgOKM5PmmPQoLkX/IDwLpsQWBBJbw4fk97y2+THK1V90oFof1AjcGA6nfgSlF8H2Fd
Rjg5zeFNgdwqU/7C72draQaJ4W7CqL+EXhA/niBGh7jPfStj7YWsj2Ou+dCfgMDYG3rHdqcImp95
yTY/wjDU3XFh2frCSHfKP+fxWRfMKSoAqsU1h9c7F1hqdb80+TnuwDIM2cVL4NX7HhYuIt0bf/aI
xYfimejvP8aeQL/XFSZ3AMX8GpwQSmIXuUig6Rx3NvyecHmtu34jrT41MtAnwEu39fZQsJHQWuIz
BucKOM4S/SFftC8NcNhTm2IHvgta3iw62dJfxSoPAOfKKEDm+EPt2FfQU6ezytdURrcjx+ltl1Kl
+sOtqcVfDSDhORDFXInGIATZtPhH9HdMmFB+a5kDBLGP7iWE+mApXWTmpZpowiCul/lMgxuXw0NG
bM60zvdEvXIthGmUeFRQ4MxuKhqKzSLoFKmIj2JOaxqNo7167Al0jy8SXWgMTWdrFQJq48/1+PGb
cF/jFFxP8NwJCR+i2fafqb4GIkq0HR+MX084MjJei3Tc3ATBJeoi9q1AHLNOLZ24gAlvUauekwLF
XcNthN4TMnbGdcgb90huWbg3t8stKK2EhRJFPjtqh2nKT9egU4+19RsnIbUqFjr8oz0APCIrC0XH
jseW3NcMrWENn7rBDzAb757KH+Psp6d9bRYkROFKUT8cbR3qvhdmTSSkvVR3PX/l//+6Vor6l4Q7
3fyLxkyqHZyJD18tHcSU5uoHpaeZf5QzkifQWr+kp+ZbQj/CwWwWVydmVQcXgxgGAfJOaVZ9k3TN
ax9egFuIvXm9oGx0k98ef7/SBKvluNCa0IRkZp4yd8bEk/F7KBF+4cIfZfIB7ntI/TZF0eJubfkc
UnJ82V6rieYOh3CK2r2yZ4EqmQdOOnVXUlw/U28cD0PGbKURJOEJgZzbXQa64kwEzcrc8Gt8WX8g
RjADLhE4OrNwG+LZqxXLtOU+mlKcwN3g8Uoz4+E4XeKU1F1zgODDdwAvXBE+sEQO18vxxbcHN+Iv
at9LwjxGeRAj3CKAB6jBao/rKbPBU2jP1NC/mtG94emYOd7DDzlyWX0JeiL8wthbLcU7RfjrGXTd
kw90pn3lRpVmFXKUzD5zrvzeMCVQE7MFvdYAAUHKkwOpTeC/0g4F1fgSxAgPbXaUqS/O6g3ow7UJ
bZYmbVSpOqwBKWdRm5UV+CnCgYlBGAjBuA35OStAKQU3L5OtbjBswE31bkG7Fwi2kEmgS1i3d6iS
edjVbOWy6QAslyWxzLoWw6JUPJRuao2neRa19ocN17XsjdMq0K+p7jYbiK5FnuxKDMgjS30H7aox
9BOoxKZSjopdXpJsP9RhH6mQnzDqGsi2W5PPercEefxV6Z1LP3wuaygqD2FIRe4jFdMXYamBzV/Y
aJzpfQSIgbPyejjjGc0z2mUQ+P/VA8mkzcIXSHXa/AXCxrPkj9ERN9wthdoA48VRA3oNl9iKRAak
yu6zUhYnrccP0VIv6oDGb4ymq5sYmQXiZqCfPVXg/S+cHXXW5GsT0LG4o7qz+T0HgFozR6vv1vGj
R1yoUb7YZEn7nXl85+wXGtNtYx0aXmfJ/9S1cMJFyJqd2JWb5btK+0Pb+18BJoSFvtANEZpXYh7M
lFIfng4j67509eo0L9xaWHich10zNvCnOZDeIH+RnbPLZQOvTUSb5KZOyDyVb5IMfiauqkg8EYNB
4b3Xv90Kpwmb4S9Ltil3Z01GloSNSdE7m6Py6WZbx5HvcKz8huFfe3iCjIU/bieGvARclUuk3dhz
cfGtgiqHV3UEbuW4edMAC3ZrneHQehRdpC/73XIsTENe7gC8ZwDi0XUa3KMAcGuF8Iy43X6Wu8hT
ITZlzno0c5Je7HCzRe4NI8Szlnl2HD36z1g0cwzxiUm8tZYfUeoQHqOc3eQac68MIenQRTvbiuAc
P1Lz3ASVP8pIs+lqH70//vWmkfIkUlMS6Bxp9k1OfLFXwEXZ8Q73aYVs1cV9FDDL2aepuegyRMKq
ihK77MwfzmP+qDzhJM0TuTXwJCR5ZxqF27vOXj8q+QKO/5qc5YHhJfx4cfuTMhxlxKpSr1m/vlcZ
c7oib/cHQLDlyugdboTlNq7V4HJnAeRyxJh2TPOrLwcJ5gDoQ+yx5M7mJCZRBAC2QbVz5OtQ4kGO
yqXKCWNfLQoLTkdJE/g+4Jxixj6m1fYVeAA4fhyop7ijW1oWvexfI2PnvsiDAxTs/ORzrYt1APkY
p0cptDEuIwMrmFzc1skrRVnPBc5jqT101+MXW1Z8ZsTJQ2fB/Kdi+gxRokJmJfDtFbmZLf+LHNtD
+FSbcyBnJIHydprUMQyOx8V36r8Ctq3alDtie4zTKQyIzGv852LxEIg89q+517urhvSx/VzTjZtN
fkF6Aradfy4UasHZk0SLjl3GLizN00Nq6L0jW8KTWxkr0Nxsl/CnZwQ8RfawMv1NM+LI7BClnng0
CmrTNOjaDdPeyPtm4Gv8+QbznYeEPqOVeyoPYpJ7tyIOueLgHJ/Wl6y0yiKmc/Ss9SKcIxzvFPeQ
yOoXgl9yZdQQFpwCzv6No6xGJfxlYEMqlfVavzWW/k721Axkh+53hHK++9g2sfL7YCiszOfpDjTm
mSslr5LuBgab6ZuwSnXmQFGOjJ/Ja0rv1RDih4p+SlqHQ353/9JX2jx4cWs6EtZK7iOZ8LK09yR9
cUJ/ttakAHjm5T1nAAkE0sW1VM/eioZ090c4KUMx0xarwDsseZefSSr+cqOI/4sNbCpx/UkrrytC
w7CkznGP8Cr+ygyCUbYAptEOYCVf1sfxWmZgR8KhywbMzpJ6TYylRpA9rHW4Ns0tMtJ7hUA6L/k8
HTOclKENY+qZh65t0ICMniJCbro5Wbt3QxNWd0v0VXtex50iL2adm8J4Dl3RJjlnOKYjRcqA1t4d
84zQXBjSzGVpnjRS75uS9eU/ZNCjSWQ06Yij69knGPMFa+iuQz4wS634df42ZjncVyd3PCYzPIjy
+VfloAp5VZnx82XaMa4RKZe9bt50xdUU2Tz3v1tZAT2nv49FKCrS3QVqAL/6SvdVNy1aaR3eB88R
93h4b7GXjXAl6Y16ceRkdEjcwHUyuIJzQP37CGm9OBGAO426UXTSfYQn8TJDATbNFOLA+xUlkv34
LXsc7Rab4qGIDfLlKYKgVRDea4kw620/TbZ3ky53gA2s3CBU5ELmCcrnEEqHoqM4/9NMDhN9icjd
befqX9BQ8Hwyxd5ecK8gmysWc/cL9QsE6TQ8rttyKNahPtILGVk05z1pWGlG6krSLFJKqHyLjtZu
FxbJ8M+mKv3qLo2Ki2JN3fN7LSybHIVa9fxrZVM8ze6W3F+2E6NKRnYzTuR5VCz3XldSaLQBPAO3
V1ky8gj6IOK/Ye+9SuahUDMcMJwEJ3ENylPRtiZHA+3InKI0QtM1Dw9sK2wyNvPstOBXPbsLSLaU
HWNgAl/UqrfXI/LtVeWTJLnq+WAZqLhvg8AMRsAGmQ19O9W985wE1VlbIf2bZ5yFl4iZMzQ9XoQb
K/p2xtAvoh5TXk1Pcc5SNnlyZExhANI8iHi/nCVH+SPICthwtQLHS1Ku0BNyJ0kQAbDJYFpsWEoM
mJKjYOSPOk72Ht4Fup88cGeAmZuyBiaQ4evQEUj8aO6Ec+Tk2H5BU/r4fPxVSjrqWqJ27W9pcH18
Ga8kdxjT4rhiqp8GOOCCzLYL2deN+mojFoaelEtmnGiSDcUdmZ/jGrmqFAuc+niZpJ23ZZ9oM4xO
fmEqw1DTtkhss1C+rItta/poEApTloFdXEa17uRlB26tp7HgverEYt1Qri2iSJQ0yhFP2FS3rnqa
UbIXvq32rJQ00d4sy/lCEUQTA5XHoJ/7Jpwp90jixVm01m6FOkswwnLP142tuYgYc4+rFtCzXlyI
+20DybUzIFZbJXKAdQlK6o+DEPLK+zjdBWk1S/HwI/jUMRUU9zrTlzm+hxpXKaJD0qXZFqhyjNjz
RLLUwCqf2LcEvd37hpYB1utWNNQWlT6VrGWxc0lMMFDgMR74iupU3ALTDoTkA3+n3/YGk0W9KFvj
F2Lyu3QLwvrn4NTuVVFlI/DxyRTNOIqmMqExnEpGx7GZXnzheFSlcF32U5cIqUsWG27kXTwUhqAF
vOCrV3MohMqP5mOyu73aiQzllnamIcv35q2T06ffA+g5gVuMp7eUI/QgAVfyivUrLFZBNG0RdOk3
4QW2ZYIQJG2VpzAKpJtl2tK1erG97yexfUZaLZ/zyIoqMi3ebtAPAMpPzPbs8zA4b271qWr/E9d3
zxncKhKt22QLbpKr2zIBAAxXwLTar1yZa5pSkDmhMesuHJeiDuIoAXkH3kQSig0JKZCEcZu/0HF5
jBgJ3JV338wyezj/l8GbQztnEdyPCizSLBsMNSzkkIyxgG3XESMKGp2OtJ2B7ZfAlJ+NYmN4ce8b
2glUWFayfR/LNkglB+KzrzDDA1iM6iCaNceDX9sHIIINSi7AVWCPSUWAeJ/+HVgESslaRUnxszyQ
3lCjSkizahnDFOz++MdGwrzZRS4DUpfsIBJpczJl2M6oP4VlVQVTwic7zulsjUDhzn/KpU71oj2N
TGGRQgxtJdvSDTRYUz/70mpIdRLz4uWwnljNMABzyeMzCBAU2guOAwEeFrICsSuIP1p8lmExVPzd
3OiW5g6W2IKg1sQSiSA1gxbEILF+BJJnkFcslgyg4A5pAA/LNPNpUFtiuysrRtEJC0v+jJ0kNyPi
Kn6kd2ONuk2rPdwgkE7mh85JuBVbEHrFdUci7oZTLEzlkvHjTbp3pQNIJD86Mgd7m30U1WuqdXUv
/JMqqMjFTOShlNm6a9VQxiLMVdWJgv5xw4SBT56GVeW+ZbmdqzCtUKgJAUHdqABGW23deE0ZQSt/
lPvPGCLnd20O13WgbIZcqT0QJIihX4AY0qGvcQfOFckKJ0dvkNxWq/NhppbLkxtetwh4KK9kHuf5
BHsTlZDwVy1WJ2qxFYoqzRMusrhI+Q4t78ILxw81cAO6gTjyayU3jGeG1yKJs7he1ABJ0QK4heBD
ooMzKXbqNVcgsIbEZu4wR6J0SeBSpazG/WGzlbTU+MsuCtsy1rapJEoKIuoAP7hmTBEWpmDsTKqD
oxoxJPkexVp3QN1Qwrrb/U9CYdB98V48eupVaMPTXKWBTRh2V6juOPm0NtbVw+V63oby2OedhyHg
VefVm0IgeuM7X+U7FaRyppgKfdL7jDFrWoRXH5A20QsFvC9r/Z8j2frTFVEFtpMNgdQXATusIsw0
X6+iwVmcrI+eezab4Jl57fUk2jGXw1XVgGh3xS0GKGu8hKViJMRHHv39kbEHTrD8eTYovSo/TYha
iR9HjJ0K+rpgyk5WK1AQw/wHrgaHnK+XBNwliv+9J6+7qcfYlbqSDGFgsKVn5wfZ9K4sG09PRGwb
/pgwF4qNZgRJrmLBSS/o1kf8bJQVkJ99iYN0uDGDBPBp1EFwbcNcqhieGt4cLfKsPRmOPYwNCoE8
7d3r/P09Dza3p/uSrRhHjozgru53MClO9lIqmPjVQS17EtYUBplrF1PJWMBrjmCYwDotXiXH0/kN
/ZECMPTmATFaav3nHmFRXOLB1GiHv3uRw36yh/77frG9u4LZtB+liOhUzJVHzUG3Hfrpj7fGCucU
eUTAe3tYmUys1HXNZ0PUVyA+PnVkIpaTBHj9LqvWZPaxWy1CpD/qdxCycXSWWs9t9xz6SU9jojxl
kWrsuKlUwoEe7c3NnPno697sMdlMRzZTxh0rmYtKT+1vERot9vqygu1uipYsaBG0OCXW1yBJI/mR
1qVnMVsXooLV4rOPmZYPmiDdw0loxJLErmrCAw+j4kHRJuvDbx74xZyllMxDttqeTtpgKxcD1zgS
k/sMV+5wYp4FnKESMRq9JRoCVWWeCTqtFXJHc1Vmu1Z2OxOKMCXiX1O/ergRZs4uxucH0o6xV65r
XA6KhLWMPJMLEealj0CEBa+6O8/Ll2SCMB5x9B67Vhx2brz/JnNXb21JE0dNQBCtYEw0N7S572fW
PI3HZnx4aeRCg4U2bVybLL+IesGq8yIpXOkchNLh/Nw8a3Yxri98klf+l4vlIRxRFhrZy0Ipuubw
1qX+Us9f7t8mq8dz178ym0yE3CMPYel9LNiLhA48B1J1hle6EGMKapQAua2oqeFgtXuChINbaAfr
iLiGspeiBjZkNJsAe4yeR8+OVOWwvtE2/HKvVV5u9RTvK2seSocxbMNj3jFOwacSP1sEQxoSwJmA
LTggOkPchqKfRRpTp2shr9ehEV7UxUsITMW4tRJ2HeJu+yT8+kmObwLhFT7tVxYqgQ8EGLCg50p5
y6CNCoPfB5muTvEbLmZ4mYymd476KKfDP+GYa5V8eceLY8kOcnojYlux3CmZOYvirAUm9q05ZSBB
YuiAn/XEyeD1n6TK0r9V+fMT1TDBOHJWEdMtamtrdKLV4YKjNQqFdK/V/ugVM3TKHu8bRGQYvHS3
xQvVnhGbHzDv8WidmvoKda1glJciuALfC4aIOdHFPNflIhOrIR6bDgA3c22VFVz6Efo6Q1JbE9TA
U8uAnaxtgmhm/Lz22CpzjUKhTpfQ8zon+8rBwxRxeY5dWeWFoHmNdd7mKk5j2C8WBMR0pvGU8knB
Go3NyweZfCwHwubjjTV4N/EE7MTtLePD5esWjcTGu36jL8Kpk/CQwcNFC1YbJ3s3R2stQ8khwi8S
SpqE1pCAmMyoC8qGo1zuckYNNxPzMfFypSAvvLAJ5VEw7Wi848eSyPAGzhguHzWf9WLrZhHhPVf4
VqqmxioqDIMiy8IthLy+PqP1kaL0vVpKBgIE0t9vrF8K7z2r0Q6H5MuQB39xiPETB/UFeUh2ucaQ
//4DdDJzxzU2lU9rO1Oi8nVHa2ChZpV4mSyDrvPNL0OENVJIpuL5Dc8ffaaj3j7v486pcLk07r3a
uVk4utAIGJGKyudduyzhkXY6WSZj78MJII7qUyC3es5kkFojy1iBfgrrlQR0NW6WEdwMI9nJKms8
2ix8oVjIG/mGtgnEjjSPeECy3FutpaHpo6x9/ue8DfAyn8ZKBPV2BtOvQPCedlYhSP5XG+djM/Mf
/NVriZNY4/6DYT1Na5k5jd+nsD2bJEs2LOHD/1X2yNZhkPNtwg86OP465OP4phBKtvoaXIYAzU4s
hVFNMYHWyCXsdngoZ5BlIwHNoQsqroI0jx354Rt9VteHBblNbqwigP5AksrcdC8UiK9/G6th/G//
vF/oMIJbna8nBqrUMLlc4eBRfGGsEBNBLwbN6wx4V/Ef2WRCZb3cH/f4Bk+vVOHLJb60JywQn/rr
Ye6AblA8+bjnJaJfB9dPbga20e7i6LGJFq7O0BcpuUYt7BbdPI/VynVzNx8U9+Ffq/3OSnUWXFA6
oOC13VD8oz2oTKUJ4PzUvsuwxMZCn4aANA0Nn04X05oRosUUFKT/a6KsjaDlmEAwIPhMbgjhpq2a
oF5LVbenmT8jDm/SHjjTOrrm/vnrkeWcEvkkGvGm1HZTODF4hGgfxoeQwUHDbB/1HjhTxrpKskYh
20+hQflSqkOGQt9p8P1qqZm54hOe/wgz+vgJ4VH6Ww6Tjebr2TCp0LUQK/F5TCiFFcB4a9yam2m9
Oea4AFP6TVYvIA7ThaEUG4q8zb/601yM35Dccg2HFukiEd11Q1e1MvK0qQdCwxNhXPrvPV8iE2ai
XDwduIQSvWx7S/EqcFPAai656KQ9i1jXODT5Jxv1FSwD8HhKoUbCD8xfG3OlFfMnoNK6UPUT8i2O
6vhQR0rWwsWHMH8Mbm5u25wG7ZJvZrdPBzXgKO6TYsDwRNNKbHVbB4bjc7taKerxSUPNSh77nanG
QhdptcHwxxuEauxXBuLacPi9fovA3YLbEphRCUb5+eaFxAKlzzqfCKpv04ZnaPeK2oLBerokxbPh
7IvmY9lc0N4+IqYJJWit7Nzavi8d0fqDDzFRBTPq7WtyU1Our2fSq48dH9JM9mvAZgWSZO1vzBlq
dJ1LQbM6s3fqfpiO5AGV9mw5+YYUSHeLYthJ8gCPzSVcXDoMgX0GvIKw6bAotSax344QzU2HfWMo
Ljo+KGlHYuzzm82JWOeJDLQ3J2LZPRV8wXwryLNu3cnnoPMYeaaNRySp68k6Vmk0ma16+2df/t0Z
YaTfWX3Z0hZv9E2neeUvfFDOFLWvbA/Yd3Wpdo69uh/CdrwAi3QST0X1GuHJKofhgXQPQxMPkFvY
iUY7zXnl3Ti4dUL4WycHdGPlJoWXRhyU9FSaH3SxQzr55t+ucWKruIkjsYxdwxONYd26xRJM88A6
k5Y4aDbjOhMl10Uh+/BPZEXtknbfMPB3fCekka4lG9aLB+tnt7L22FOPRABYfmmWAI4GPABt/ZSX
gkHdkv+Qg1AgXLyANWqHTs5pnPr2QkT6JHoZ4rW2GDYn6aIbWBnustUfdjsBKTxtQ2wKd0/idGUR
Df68f01o6tFihGAVC3E+cRmFQluiQkOCty9COdCKxZ31sd8TCXHAYrj8XI1UBIqWALRO4f+7SQmH
Bs84y/GfFwijhjEFTitddFe6PGFp0KndY0chuafmQSsvVpdyPD78VEwISNi/sF/1wrMzQQol0RAA
RAgAwyDUwmjv7rzOd76Vy4cEEpZb0t6vS4Peb8Y5fI5RVs+Vb2B6LCrU/W9/sRSywIxJZP6CdHj/
hXJwpGo3JXAPqcFAtPKAHI3PlrLsant69Vg1dqJlK9VU+WhpJcJ1JTFhx5gwxEO02LiGBmK74Qd3
DhxhV9nRggmc6THZYvksfocwqVg+V0BHlQhMDPIwd5tIEWTqHngwQ3n58BL599pXPw044fqEPrx4
eLTL4PWXg1t2g6XQ9IFfm8CnTairgmc2+DhTB8+MJFpA9bhLOGd7JDiI2aTFAWX/ZZkw3k9PvlW/
r9oELkfRdPl3WqCyT+1DEKvQZbwL3DXWeABGYColMz92LuuzCsLvbTVclsReB39LsHELx5o8vKTr
X89fDU6vaXM67fO7o5UcHINn8eXMpIx6jKt2CQ3QybMfjVXjHbkjyrElyJJc8DjcBQYuS63u2Tt9
EIhpVefyPppLK25+OBgrypO7ZZnLXtN5Z4SDziMzPsKJII97vs8B2MK+v5b4pCjTFru6MaZRvATL
6AdXMtbpu/awyT0gpSEWopedmokH2JvlghazGyA3Hoh/4EfNLlh/qnbeVTRDShqFg5ozsM+aiz1S
/KjgDNfDZZR45ajziZo5OZYmKHlMGPJ9QN1jSgRVE2HPztaL3nyQt0FPCZ35b4svKky77Z/ZJhc6
FJCXeBYL0K8DKl052aLyeBxTf64AFn7PWpBOyxNjrR0VAqE10EsVePVTdr6ar3yGxcD4aMvGEy/L
b2dBESZEg6lZzhZvywYTzTM1Atfpa3PGW0R0HMZHlnFgmeFq4fV6XKAL4kbVH9zmXRyYFONavYop
Dp4K31qCMJvfoBvzO9whxtZgVfEAHHVqGpw7SbIrfLO8XswR53X3p1cCIuLD0O4S0kprCNO6Z/Ev
JJkL3L4k2Jtc2m3v8iQiYz6vwQzhl+jvyv0M5VB/Mpwc4J9NOx6lwlph9Z3M8AP3Z2LiPVn8cvCp
zfhxrTE25p6dNXhZBiJP/8Xr54ryCwHtsGC9xarK0n9lviva2PDnJIUUVZpsV9MYOA1vDOITXwsi
iwnxla1scZMOIx9/GeIw7EEDWu9VJ08eE1X/KdAgE8SHgnAeeq+cXfQ2bB/qI7fbcpsY8K+7EKzi
rD6/G42lg/L//i4fldSaJNMiKJ+kNVfNorZ7mMnfG2aZ81bT27pGe65glyxEGA2fQo7hv7nKUHSE
5vm2MZ/wBdbcatcXmJujcVt5eJb4LMbbFnR+CiEJMVZyyOVgRtdCs0YQ/qbTVEV32Ap9v62nzw2D
c9DU/Tj0uUQrVFTuLeNW9rd+o19G2RySpgVWQBaxEwZevgG7VkYdM5VcS8ImRV6r5fWdREVFtthb
SgfTtHh2fqKH2kf8449bLe+lsDBZ0utGVcn9yvGbH/IXML1xi8wUHRIidxw0nzWk17LA7jIrOR+L
Z75RN7XzQUHVc0kn03aIFMtgwB7bUwNth7Kw2TRqBNizip8qtQ7fvjg0ynbmnfBM+3dYiYp0k50q
3hi1EyQtshnY0h6jdBgf/GsliBFtgz/ojLASNtY/fLggwJWDjktOV5IlpZ2mjWHDbBmP843TnkXC
WZbE+2DwhaaMdyWmPVtjJfnomoEWpvmmLne00cN4roLCGBqAkb6dIWXaOiqp/C17d0CWzaA6U1M8
GP4ipoOIlXEM3HdeZqO/vw1B5nM/9lUwU7FZ4sJEMzdb56lblygAEYL9h0MmrbUjbxRBysdgnSPh
OKoFvXBC2IvCV++4NwKMbwpMcuJTysOM6GDvaFWZfism5MxFBW2mjeYgD4i093JAjGFawmpE86pr
DK/MyAaZEgJjTZSWKRU40SXW3Qd3fBLqryvCxstJQ8YE7oKZKlmAyNTvJYMipsOoteJiTl1o1/P6
KhCtyGPWiUhPHcTPM7xDj8L/yOjtqZac1Wtkf7nzK4EvPkaOvMG55z6cDwj3/kN2bHILbF1IitYd
gNKBzxnyOGpCv9f8Aqr1d0O5htG7hqSr7sbRwnj6TafT1RshWc1Tx0pF87aMevRMpLKoKS74F8Px
GjNox3WsuqVPEiemLKxYz3lyte/14BXbyODGEyR0Gb13Dp6NUbvFP2Hb/GTq/bJ1ChBwcCUhzMAn
DFYmI/O1bzkHgObUFnbOAucXRS7BsOmgSjBr3WF7GMIvnhd/lI1hdIOjNDG/JmhaASvKQv9uwoRI
HSR2C8RAmqWNWcDZje52qR/t/osgg9X0VeAxIwmF8i9eyN/7Yi43/bptn+QYREMLOd/oKhNQ33YU
BOmlY5qBizpmo7bONhLeBcmBqpGyrvR+RX4sBL9KhUim69CVV7V2fZ8XuKu8A+uy6wZJ/amFK0vI
5zJ5iZ7k/NVazzny5vrHbPKgfMG6MGiwTRf1aefOhJHs2wELjLkFRiLHZVaSkP9kycmae1PcmR9V
UEZQ3U+hA6jQfZAIcX7Iq+IYVBuuajsz00TVXF3F+MAYTkyugNAUUrYDTNOrgApWeQKvR3f3/qDW
UjGwMFcxfugPcMNFueLYsAlD3RBCPGECxJ4Pn75R/sgEm+nORk52AxwF1c2VRqQdrh3aBAI59hoX
lVw2girMw3yoKF4RIVR39KeQ3guAUs7uHsDEB0gfLPguxcAggXVGFNDib6cBtr9HUlWk26L6+1Ub
AaJnnPMfm5fiSMQ7GSuIMk5xmVXLJ111Cswjb356hX3broJdLVqzEuvQE2lljzI1+N5p445LXYii
Se5pgg9VvrCnNsJSW3NgoxdBAB6dUckI8z4bwJCDh0I8oqHhzB3699H9uHaGLlWQMO82S5Ht7pXl
0FbQbROd5sNNzxXaL34huhK9khunR9C8UUd3o6wSeIN2IP4PMH8CJdc0shGkXBWPHueYCr1o1dR7
HvTAqTRHpuPSKaaAU8jSsLIq6RNZ5Wirg4a6fwnMPirxtbeic0F/VNbxxSfnUmuup1jPlCb0TWiz
d8qcMboXLsVtABbcIXDKY+BOR7gmy0l6zv2eJjC2zo8X8SJlDixx5IAhWp/HIznFn29Nve1jgmb3
wRoZtY1hJt9/g96WcVybjbyZHTp8in7Kmg8IS+RbZWFgTM0K9IV0x0N/utuHGc169KjmpyPAC4cX
4ICNls5FOT9Iud6KtfdGGE3Ti+DYrQ1+N1oPZfMgjx8wra6w7XSHrMUB87BrQ9nFivKdqsWFt/sT
1jOAzKmUZ5Jd6nz9MeybjQFz5Pa+28T5XTbXGLcDuP7fxxgDV+wTzbNp6p/IU4RBVn4u6YL7xLBT
QwnidU9AkgmtWHe/iRowVc08IvQDba7089ZbdSNMSvLejYE9kjn20PGjRwrW6oACZZNsQd7HftFi
lptn93z2DZh7j8ajBuwIPT6MmmtingMXmSx4nbbJ7dbR47LTCsjfdFhA3OGzd6twgo7XtNOu/L8n
lIIU2Ka1Pr9Qh5V+OKEL5D6LwWId9H5bUS2auoXvYWnhZrJh/YMK5JVlnERfBvT1gHszw5FC3NeL
TKmGlyg4/mGOGcX2Ayk8UcBb2wpSyTwnjfwBkvB4YGpgmoUfmvLL8UDI89oUxGRL0PikebO/z8y+
f9c6lNiqDKslrLsMnnw+8TeNxkRrnp0fSdsL2433Ser9TCCdh04GQQpJKikUUrmySJiV2nRpKoSV
xAZxiKysoAbELyn76cB+euccmgh8wbdJNNjc8b1HGTzkSu/3D2tiXaaz/SZdTqMf1mmo3XaiT7Dw
/MlN7nxPPGD5iwreir0SH/v+NbWh6qapzylAsYq7SiLbmW0R4wKEL7sJ3yRPQCzQhVpjqpGhDCfQ
FX8iLe00jWI4a/44wuPITZi+TRVkdmBvkIxtUSeiwj+bg5eNlomCTuQfN+e2GW/QhdNxpJQiKsqa
wPhgSiDoMUVc507Lg2xBMaeygBqlVDo3tYME9hyi3nuvI3Wz2c6MQvz6+BjtWczxlR0q3tUr3tRx
AMQLH/ewP5M5RXrnqni4h7DSKeDrS3FEdStmuI5IDSYabIfQvUAGaFUrIQnmWdMS5yS9/sGyqD9y
kqmTV2GafmRcnjzBVOxrV1wO/fAoxWFyKGm8I3mvYAMnGquJUNIlQL8y68BowdWf9uXijU6QGBqU
N0jWxv6SshFTSiGkuDA2y4noC02TmehDj5U1Yi1B0xXq/uk9sLN6UoSM9SuroNamDalr7Ucjq9is
2UtPV63HfRIMdpMVKTLp2Pua3K16vrtRM0kLcoCCX3zpdHkHjspzpeCUOV6Bk+6XCxIHy647vl/v
TLYTfd4ZXobI3Op5Zoy9kkhx4MCjRuDc+l+ZxzL+zOlceHv00JzJm9jnm/jbl2kubIBLgxkxhlbZ
6a2OYQW1oEwS/kyH/sp/QTzASDLlS92VO6N60O5wN6O71TRe0c6Vj/IKwo/funqetc9jQPtzdImM
uRFp2Uy28U2UMFIyANpO3Kbz9J8i5Max13a8N44alvbiAvGnAGqmC1EU8LEwhtKSUB3gD05L3sdb
QCnscNsGTqVxZ3ZOfjDoRYFL4Jpqj0sNFx70rn87Tjxs+DwFsLR3sn0VxJyi5aZwz314naNjq7Lp
jfTaQ6omBoeMYatj7RSvR8LrdKU2KmE29qfSkKCegYRaqAtONALAldEL44XJEaYLq8c4EaUxg7YT
/rcRI0ubO7zihVJz2Ku6y+xEA2TUOdruNTy8BcajWzQlhIORkN/fhDvJ6wUoXv80FbxTUJXypy+G
zznoiyejeQLzEcN346xEgVMqKaAp50Um9CZjkjwpTle0GF4oIax0kebjurze+RxXBabkd3x2zOMA
1cKY/4X3MhogxrH9j9B9Ezn3FT/WivLom7p//69jySWTIpdB+wh1IMR45IVHB6Ny84MIzPJvQ499
2Ofhr65CbbuIsrDDgue3+8iJTujf+n+jqvOhPiczSP22x21zaqazkZjnQ2D76PfcuPHB/2Em0Cnd
SOUNO68RrTwockmblTtPINCDBnxlDFMp4MNFiyyiKvc3OunEMW6q47SvzqnyfgFYj6mtTvV7nfbf
wXMmHXZ57vf3Lm8BkkbxwB258JWxiro/tcb/kjTg/oIbXqnsAZCk6PBjkVzNeiGDF6SCvaKQX11G
z/L7HzOYftPodHlWZO1FJlMSMdxeF1bS3/JSw3SEGH2rbYh6aOI3hiEttTqQJS3io3Xd8+7vrHiL
NWrUGgTM1uXWFxMaKAMEKQpGRrfT8T16j28JT+qj1ACUEKulT37bSk7pqhQsZrBibMNWpy2ZB0Ne
DrwSkdRFl59i4jupOgDUL98ieWQGZhfZ6sdcQIbMo4QAW6QY3/2GszOLGWmyfbjF5eSVXpK5fPuH
OoUi3vX2uGUWLbfaY8OGwdaxSTBQ4OgFkshu1DgczxduBQ/YpXddEJy+My37YQFrizOqYk2h6qvM
18Lu3GZXAb1182yHt6FNjDbz6MnbvsRm0Th0dqYYjzb3yimjg67FJg6lZIPRc+JQ+TCx95kR5Ny4
ogVDiRnjnIo4a7vVaPrjyG7gyCav7wivAA175R2z+y8YmcOkUcO1W1/KehLR31sDSmKd35uu50Gs
Dfv8mtyrVbUlSMFZ+i7VMll+rC9LOl9YLjYgWlHEDq5GATm3Uawcs1q710sY1BxySzs8EQjBM/fv
3TqNVAB0WPzBGINwgpm4tjP+l74yfnCE27XFcxkOOZDG7f3EoMPm4sTlUdoumLcvt7O5+DyNXt1B
cLhNgIk6Bdpayq8o+9M4ak16uHoA5p4jPzp2o2PJFT3zFrgxd6ZF0NZi5OZ1AMoAZ9aqb/nwJ1Z2
F7IDiIpaD3zjtaspJpt+sfyun7nRh1LYgqkEJBTY5OyODxMzcIeQDWliEEmYlgVhiOKJrJ/A4Iri
22Hv469Yd9m0lblbhd88j9SD/qfjOa0aTNJTtuO3ZN63NFYxCS/FGSaa6LHYvK4WCYFTH2q39k10
uWm85RWfv81D3tOk5xruRIdALnZUks9hsG5oVnVJ2NZG/3sz3T1SkSBDmDhYzT0gczsyex4aBZAj
2LmaewROOkXrbeqmT4CgiMb2LRyILTjeIoBYCy6RGLCRLH7gJJfIlpV539G877cahrw/LseVqV5R
dEAb4bVjknSQQ4e0IZEm+HhCT6PQvxt7avPF/mJmyypmXEssUBB+aTX8AaG/AndwK1q0KQ6hB62n
qozXE8a7IU+sRXi7X3P2PwUPlS/2HW3n9gLDbco/ZD11Xh/5JuVBRKFxoOM1aY5r7TDZxvb+eFgD
TM1d8k7XtvWeRJwWtT08M+3aelNIdnqE+3nAug9S9cWGbU3Ks1hLyY4QBKNlprCGqV00j0XaViyw
qLMQCo6KG+sFTMm/MKJDa5zpitoMFrOJJRcmNRxUnnh7H+0Ie0418EVLagEWxf0nYq1KcCUbubIb
6TN/c3j9to8ZK3npVLzBJsdWz7so+tBv2vfIbCCaa8jXFDWms7x5M3MigQroY4GShcD3jFE+fY21
DuYxTc3Aby7C2XDsWd1m/8SddG89/6Yrn5Vf4rbf9vE5S8X7ymMaAQ9Mj48YnCs5hgRSgZV3EfUC
fgwktyAfuCpLvnWxhSVS12T5td77s+81d36hqc8j8Lvo8zVUTpjC20WZsD8xpQPoaUhGqJSWsbvW
Y2N6NmvGZ2McZsY9z+HQPivlIi5sPvV3j9a8vX3DbJnxGsitvluLWb4yUkgvzLRBRBaW89/NE8tK
4acTYc5lC9Ci4qvwSUGXo7h8sTCOCChVgVHH5D88gEHotGkiJtrRnfQB9lzL8BhyW1P32jIl/6ZN
d9lBtdl42//O4MOkvmDHtp9NIYK0UdsEgYok4F9I4ig+DJ7F5pwd38RVoBHIMVRxOtLfotbyJK/E
raNzMyQpraVd2ityKDlxB1DqxUdZ7pkjH4o7ZIZvjjOeJq9CFFHyJxEsUgzRMszhqIhaHnHdDilX
gMlAXcs0HROrnNaD2JCNB/pha566Dfeaj8feUPw5o61W10ITehoy5CSM5s9zwVDizUtgsG8V9B6V
W7eqw+hfD3QQgS9+Y/4+xP1z5jxaJiQ9rDonXOBdoayYPGS1hwpoeturBYKJaQQo1O5cDuAio6ah
R4KExyJD+g0ldYqcWJE06cNV7Jw+dlVH5UXbXecIbVkhH5nHeZJ7Se3L2PTLr2ks33X7Wf9qI9bN
SaYLANEzSo/sUDf7Dvq2pCTb+0XkqX1JfDpNWtoGM7eb2B2ALQ723/PQKKQV9De42GnqL65LNnVf
70W4jYTyx8PhP7kiG/d7SAJG0WtUV5uayw+QyEa7LUABl2z/2fDtht59emaV4nwDVKcexzd9ZYaP
9qkP49aEiZndNiNFLmtRHUwTRlb1ZpgcitKItv3alyiQ7WrYzeIt4zmODYqyqVeqJK261wdEnuiB
nRPxKR9UiWJ4GJwT2Mk6CWjxO+VSroV91BBjbkocqMff8jpX9IXJISAVqDTzxfkrAhxpHDfoItTs
K72zo85WnJN5xPxzlxCPX19Ji4q8qn1VRBEulrrYD+/ReLihj7vtGqTMyYke66pPvWBuNYvJ7eV+
ZgT2PEJSYaTYGNXIX/x/erJIALLBC/mtR/1DqMuK9eNGZhsfdK04yIYLjWnFpFNiDOfbiTWqTJC9
7BXTWrO5eEPXEzkSluPTKBRv1Zd+mIZy84lk/ttFUJSksqoSXTMYVmkvmLst1KoyUfkU9EGQVR4x
uOnt5Dy54pz3A++Fd1pP5v4JNKfU94BQ6TfJyJxaiulPsY3w7wO1xqtYR6nhiEO5st5LLArBiMbs
xPFTa8RBlBRPanf1WBq8hjGPzR1Ito2sCQjuqtP84lT84OXKEiwQIYdvwTbvS3gtDJhGc9fmSeGN
LWEKutCATy7gAPk5R0Yud4kQJVPGfic8DQ2p908b25RV9dqDW7O+pv7YgyZ//GS496W3wWbtmFr1
RvGDrjy8vmYXOvE/MdDbRvhEqmDn/XHBNA5DXeos+bTU3UpzDD74f7gwid2VLuYpeJD9dzR7n/tS
oSC9yYblm5UvEuwWWJ1qUG5KynmL4PSL0i/egmZd823uGl5D7fEA93QFtUHqtxFn++NzzbiJK3yo
gN9vmNrWCn7W+VtnKUBEIcLRwyEA6cPFqhn3E4ZCVg6oYoYZNt04nP5RmXp1JGnj52V/tdb7Kn3d
VYJI4XOrkk0jyDmUqjoFcL3CLHmhapCPhLWTTTfxJt4xAto4uMBodl88ivDQLhV47WlnXtr74eHE
sbd3NBM19uavs+xEnQXqm+6j4x0dRehsO6on/Wt3uv7X0dHZ2uM3hAgX1G2eD1LFsYP2WkI4eaMV
8FrT62MQ3f+iklhnni+hI8zPYO361rkMt54IrcB8iBYbX0Lm1u094gMcOxvcrPZjWP+GhzjZbJyo
OvLKg+pu4r4t9fVRooaZmSRkXmwWLJS0ES/PSVci6MN1fehwU8AiSjOE6uAR61taVn2nGGot1/qM
HflspZkQpafyCE3g0xfiapXbTSjSbkmcllc+MkjuHmybup8z/CCHBZF3imhEHgxdmeOdKU25b01N
KrjCzvS3v0oLWaRcit/W41ht96kYgWh9o08iKr52eZfIkYO1cytGcBr/BpSjsGdddQxEJz9TtyAJ
HvZC/P/Vhk9wh48nPqXrFpnunjUDr2l9f1cHRMbJjaTUVLGDnkG1ZpNCcVnVhp14PtOKjWM8vmHo
smTkObtdCXy3NfPQkOuAB0KQ1tAeUb4e/rPESXeCbNNMaB53MqUorTumGuoVvkYWnSJ62pj3u7Ik
VOU2XJONoAHsi1aJA77iueUnecv1rUwXPJernAFnQlUP2UfEv0Zoql2nE/tLFxdjvD527+OQiBaV
sSlOUqtrgndOX9LuT8iE3xmYRFz35jVXqpZBDCFqVZhYXxpuba4fi2DZHRf5obe6Z+JtKy0eiwlY
zhLJr3NVTpNvquSz8byh6BdiG97eyuny01L/z1O4quJ298IchwglJLW1rgk5BjV31ktEbG8m7kHc
A3fvtstBPGX/OPUsRsCvcY5Th1kYjb5sUU7gDFC+yuoeImRvXiEji8kXbz5DDtt5YFy51WSkyqnK
2VYxcTUg0ZvZUZ0sDXJzdtckTB4ZikBJ/xt06hDpOjSEn/4WF3DJb61Ax/LYsACfjzVEJAo4NUHN
t1lr/PghsgWvEzlsVxvRIFLQjvuSESf0fWSwOjrYLyl0TWyDsrDe7RG5XRrDW0pyE6cXi58AY1zP
tKCUK+da07MVm8qaFMRZDugD8wYhL/CRKsMu0RWb8BlmoHji2S0FjCm2QnRBsWlHSuWPnPYbOJlq
q8EMAQ+7E43ddHbx/kVqgGMUPcBgEgZNlKyeoAFNzeTl+g1/fVQxMyLdPkuSDS69UfWHpUl+1Wmj
nJUSWabU/4krfNLpzHmBltXkTKHpH5gRXRPTUBwOtl31gIkqhStw7o+WY0F4C3ZrDfBugcS6p4aL
X42JugHvUKsNXiR3irhzRt7WkK9sPh9VE4jDN/mjE9ckTgD1P+FJpRLlkejSSr90PIt9kUn+NyW9
J/8YYM2w5DvENmQeRTt4z8Qec4WSR8aCuce3+qQ29Z4/U+nzwoSok6LprM/crHJR0pKpaObBX1NY
gNs7u6Jx247aXpA+lpfAFZaenV66cZbpUHxKyxX6+6IpHzSvI24ivggnHjHxFDhLKJGXpxTAL3SC
8d3uF6sYDqEp26I7gl6x1gM2soyNVzq4umw4K2ykYva7g1QQqZ3NrtmLo+izJPkaUijLD7H6WUaT
5r0G3LoBW26ilShALxlqPevbK+qZ6shM8NCxOOXEnKu9Pp6mM+tjQGDK3fqGBhR4foQXsSleEZUt
Ddd+N3PhqmhECrbjPxaWyO4ejwhb4rTATunsn4mXaC1BqCNq8nHBZrWBzS0sE54B9IGarQ+NyqrG
Wx9xRbNCqcbfHHpJWd2BqBNSXOXziL2FJSk2yR6AHIVeTAORU6DW3LXxN/l12k8/oqe9+DC5LIkq
MiELk3CwZYJOJ3joYxPap+1p1juwjVPbnO2DGz0C7a2tkAS8ByRS8cgVNATrZrdqJwF/KI3Y3Y9Q
QFGdmFi3eQb6pGWNljx4mDc6By+pfEv94roos3iE+KPGdWieu5SlrVMKD4TFam9QkUCX0ZSo2jja
mc6PvfzdjhXvfVMvP43IL92DtKdvbRzmz8WW8tH7d9fxZD0ihe93E/wrlRt1ZCWg3qcsUV19w2w8
jKzXMKnhPR/Ndk3+Wc+9XoFNDEHMaF9B7uku0btVFv39uwRKmHWzFk2XbTPRyW2qCRDwPF0vrLx+
X6W5oInL6xSRHz6z3zPL2BRuADJhGsS8d4B6MWi/sDsofCKe7Zepp7UBKrPajhFzSkxc/f/ufx03
zB+7CtrGWxObdLKSJZXXPqjwroDfrATBai8TV+KssOwCvfwk9J05Tw+sa+zmi5zg/99FMfvRBgwG
F2vMnn5cp3XZR33VsGg8NMhAVuXM2Pbr9pUb7mAoGI4iK/u02EIAx91G3nbPa49dPXvLfki54oRm
nDf5OyfJiRs+EXOktxF9Q1iNWIiD7rKMjzuTJfhhW8eELN2xjwfP7Hjk6ZTK+NRqY5zYbGkgbWw6
IHldd9CwqacrlR4EhzjEZxbh59Ybx/wHPB1WVuh+KooDnjgqi4xWGaV6pRsUALdk0L5uh5tpA6lT
rdSdQt3hL/MkADno7ELhkNIpLmq0Hh6fgH/KyfoCyKSmeCLzJ0U+YsOi2kgnAR/IPtkk9f00tlwt
9ezVdNd0qugmwnzfcnVxJoGdAOVNWn6GL4SQmgiWEBA/62w9UXgi6gfGQagkFDOaWvLo5ahtf1Ad
YhZ5fuAeJwQbwaafDmUzsdFLgMlcd23ATJBD7NngrwFgN4wx4Fpklq0MoH1fDz3mVqlUJkwgahM4
Y1Mjga98YomQBFPyyQsEpBoBzM9QEDTohW2P723n/wPnEyTHqrP6Pmbreh0Pfa/3uOhd7hgfzCKr
VZ07RJrEU/ri5irO9lZwEWSjHhOEgnFqycD9Wmz4qtDl0cOHHrUrT28IHNYZuFX4FZb7pmonuCmF
/SQ+91GfPu/TML+bci2XaSPhjue7n7GRJKl32op0+lyGJ2GhDh2AN3omCm3A1xIXSi/9TG+LPywW
TXYQThVh0W3dzBRCYjSWqXJk+t/COTrQleqCnnp3CAi3BOPNowmrOaJNrdcN9Fj2lEcXUzDzqkX5
4tiGrio2+ChLsc8h/4NPp5rVzeiAFM1uah+2YQvU9InUd+Kv+OdaEIwF1snR1pD6Gu9bYel0/QoW
KWvATB4QzM2FTvVeeQ+zao1NRldYa4QnwCteqsh1vMQOM7Or5N0XqHq3hJfQLNZ8vG5oJsez1/VQ
zp2tcL3S74wUNLLSTbofkWtLu12BVAzXnMo2Tr6W/VkLVGy6ccPQMbvJAQPci2aIK2ZUQLYGOjfg
CSbo/OhD6CLsK1hugYNf2pWdvrimceW7/bUk2oMiUA3IzHe8X7sg2qS6Yl3alkBSufUGb0MmbzgA
2uCa1bzmL7M07xLJIhWkpBM4CzUZesn/xgeNUQa1ZlCUADzbVSYesXm6N4a5gHSctYMCK8qGzwTZ
gWr7CibXhSeEK0QkJbCOAR+yBuyhBPGvdJtPorCTEYRUM2KFQomh31hpnLbcKpaPzYN0L4dYDX0B
8rNad2IhanGdy+S+U9pPUOP1ILq4yiH7k2SPVz6LBz/kliaEg2FhrDqtRGUD6zODNk5AxtSEmsXJ
oeOoYH6IQhkOzuNjKuOOX2FIU5rUvftO+QqOaVlPSTW5OEbPuomJL2LREAlJPEBoYZZNlWoVNVrr
bZtKlexrIXP5OD8vWzwpMpaqQ2ugvqS0LkoviOTO4NwqcEZ56u+AKnpvAoeg2OeLyJ7OLNNYaPOI
gwppfb0BflWPKwrO0yef+Vf/TmmvpqBr+InfiE82+k66eD8v0PsiItR5r3LYBhE0hrCOERXBO0jU
RUjqVsXug4H82ORvCMeMoXbE8Z0XMJtu+7yBRlTLYy6VUpeuPwwKOvyfHcUNH6R3258cW+ZYbatC
MAKzfyVMCLdyjwuQe3P2halNdzIZJf1GYa81uyGS9eNz1ME0+lCztHmtb1ot+g9FJOb0wxn6Aako
tcPu52D4sVfUCDmwYlrSTnoVUM1LmFIBYEvim58FRg4JuNugJ1hvFarAM2I4Ch99yldB0hY4Pn0P
GxCpf7v8sad3SokJdPYKDmK8e0gLbnKhDvprPYf3p2FEhlwno6d4IrAtWq8HHJDvZW8o7FTunMC3
6lP3od2CjiSZRsc7J9VBhmBmds1ACNnoZZG3lo8ztmmOiaswhK/iQdqgCdr3hKvBxE0USja9R9Fy
4a6C43zwrJ+QLlTVzfJ6yyt9Ucvst+FGDxpe8FFMRFC1czZKelGVsQnTZWCveGXPWPpzgGr8HC3g
vlstIll+vTmv9QBmgvGfxo0Ndae1T1voCHzRtRn4dPOKBJDCY/hYKvU9twsZZmPaMVjEoNifReZN
2RYS8qyBG/2qyvUmG0ubyDeF8mrola4jQM+jFtC+XfZ678NWfmZDbtubIjeAKHVF2B8VbAfOdq+c
OtM/puPstd9GG8gPGlSso8Xv+Ndoq9I5o+ISXdcjQKo5ux3gyyCzefnXyGVg3tOTmiWkAPBexx6i
AublSZtwmv82s6rhsFqtJQB9sG2Xdhphjfu7s6Ys8fdnGaLBcKcNIjXWMm0t/2BGOIfdrFDyTYWK
CNzWAWs2MNYwhAMMPenPIqxunldFZNn1XsZpNN5cZMS6A4XzsuNT9qWoGNkKU90hjTFIOheB4+5k
VNWKhAyWP9EGHeVtJIBn+scbIc2ENFjYVVSU2NtWwqeb8drnfp4OzOeV/2gPBppBxJsajbLwtbyV
8PSk3lKIkw8VoAaX7I2qWksX9Kd/AldB9mrlDIN+7KFZwZZJMKWQoGgOvyJUEeAw51m6poxgVT7M
SWr71qrjLRRBlryQ3swe5RTXvfeR8/c2IYMrpBSSvqT8gY5PkM8EqDEdJxkTWPAXgg2NW+bCLWpa
z8t83fEug+8xZD4NtR3S932XPpt9N8zRJA/okYDM8g6TV3cQ0yQ1Afem/35iYkPjuHXqz/XOxmyV
T0rPD0qjYKFupw7ymiucfSbPZ/2sNaG4FdHVMLfU1ADtNY1bZDvS5uiVxbWafaKWfhkJMFkEFkb9
VHnRI7CDJDKD1++qzOEOQ7pnHhS1Pxrk1b7+3su4jDOlCATv8lpifhxY523sdD8+GGm1KdIE7Exh
f+c4rlhSotue5IP2VU+kh2nfG1DkZ4095U6JN9Hbw+FrL0oFLS7dB92Z4ymqOEpQzQSTXOm1BEKh
A7Qa9xtQOMofQWbpCqjPwKpLR+S8TQw3Glzp2vYKk3Y3AdPZhDzZ1yI79qt7zEJ409N+yxcN2t6d
eDwMkKvUVxIKPD/SM4cAgswGGiGD9ic3Q+7UEvRJWIt80NMRxsM2UJqhosDzafddwMMGwoVHI50E
g1fqHEZ7hwxWn8WgescUglIDdMuO7jLVf83Fsvm4cc3OrShz6S2jmRRl8fj1j6OnuOAF990Tdw6m
OYNS/tvahQa07AivW4eLgu9nn36urP+MDKu8Y/mkoKnN36tTv16o6kFCsTT3GoDvcOiMBYsis89x
rdRhZRSVhODDnDasenE0gw/Bn4nINSbsk0zfspJjxUXrbu2YDFNgu/DtA0Hl6PExUBJhxeZM5fA0
L7dNgPi+DnrjwK/oLaiTtLhC/h2LDUrlnLb50v/s1UZyDSGFH6/FYqsReBtZ+CUUEt5KugLUb6y4
rqso5vRiN6lG1z5KFe9me7g6887dBntH+mnVMkcD3MZt9x8HvC5q/aCjbNaShhuAXU679+HQr9mC
ZVGL9ec9OLsQUIkHuuub0/Ew4knnJis4kmMz0bTs+WgAHxykT0p7nj8nF7LdqXbnnl9iuAsqvJ1V
ToSK4CUK3d+1seeakV8RRdlDRoFm0rvVLRBZmdrpFVHM/Mm2YZiOnMQIb67oUL/T60IqkvZ/ron6
o3xDM0EltlZjRF0GT1ZdE4JIFhN92wcSEuu/JNuuxWGOp4rmPn3bNYXBfrfjz5Po+U9uU3EqJ4aY
uEt+LSco7yc0k1WC2Xj9lk8uy0NAVt9qtNu/KRV9vo2XP9pgnayCtcF+nMY3uC3mcG1XqBTR740N
CA+7grM6XPKgHIJdlAOxo2F2CNALNiXzmfuuYDQrE1Pkq7TEcWStd2fln+zesBBkiwpPFDXNI+yi
jBRVX+SLkcBoWRKeh0ZQLuPiZ6wnWYQJsRyDyaJ9bVRbGdpvtO6cbtql2oVK8jGWHQx0idu7RhmO
dnea6EmZok5ksI2AHRw5e8vYT+Y3mtDwCr2V0XF/2A6A1Uxkuy5oZ5H3QXrNCSO8zPMN4z3QIRVT
SrHIg6JeHSCb2PorpCaKfDQyVVuQhSzURKIPZOEtCrImH2bPCZVlnt22jWbu8ZWuCpzk8awQd18C
hhji00Gs//ybA2l49++5DGAodngR6Q1pg2IV8cvdf+S+VX+imyOB+hAxGAr3SK8I3tLXgQkV+ybk
mofWbfgB3HQgd77kLmoeaEHP/Dv/CCZsRiIuU4gkbAZQCK8LJZA+cpci3jrKdnKcW/JzEAHjx9V4
AmOVlUJ70iC+44kHEDozI9Hn05zixDWX7fUEbNz8PgxFSryOWU4T6yWeAF/82Iv1T2rpuxzQQIln
nwekAYkYhVYakB+K69IFZSBAEIAX692319Qa7/az25Y0I5A/WSAspqZ/qDNEGe52YLHpQn1cwIaU
QcR9W/UBJv0+yUFLYe7VSg2rzeturxM18MGf6o9xmvMFoXV4ssEezU+Y5106YIas/Ar9qshQJXaI
gcrV2pXaYs8MOTbaP06ozC8MQmeczK2+W5/AJDJW5SJkGpLkdZRJaOB0FB0TqozDg886U4GXWX2i
MV+5QeD5CvHyxTBT5b1u9JkSS7M+ROAES/uPPgr0j0GwfNo+FKAWB/bX2Zpmvz1Ct8ApoQigHDe1
/rLcOUj38D+4FzhE8LJAFsqxG5wx1ILbHzORhLlP9iIKrmAbJFY51FadNdaWKjH4dQUodrBj4q/1
b3U22R2YpbwoEJlc2cr5gpUIrGdjZ2QOcqQ18zvi8kkQon7sRT461hMvwXYAp8EatzUZqlXixNTh
9cwHuf+M+2Wkku1luVgD4rSvRLaKD3HWx5FN5p1oGXMjOaACHqN/priNUpMwvUjhbSI4LjU7RR3u
vtWBQZ8nT46x3MvzziRASKVHnQs8IxSJtH3Ltd/eVoy4EsVuAny/gg7sBN8MIPO+mLkz/XivvGer
EivpEl95uP3f23tqxVjdNCAyxleid8OB0ARAodRmUHIVyz3T9n9fOoleC9/NlslTkFMTJNZ3X6MH
fCIJzmjS5ybBXRtjyNIKiUOlVSXNJrTAGawtLIFe9KYwJ5FZgkr2Ejq3pwS8ol13WYHcGAGQyfFs
731dcmpyM70Nyjict1VYJGM6HPu4aB4vntuT+q3U9mOy4rhYVXQwxwcgEDpi+exfFFH/wFEfIoJO
18J9PLAWXQOVE5W7r0PllFUzhiYkJ0YaDNDnphjdNNPBfzWWKhn0q7TlUuwBbCEzbtklggNeuGjm
4+cVLaIFZOlHt769Du0nFpOx20Ee8pA9LCQ492umbNJQ/vwz/BMr53HmYReL1kELR7/L2OzgzPHi
xM/Y0H1UohkNBWBghYRDez+5sBa7J+a509346Fuq2dgGZo4o5mu1/iTSZG5mzStCtqQ1tjGdkj9y
43NK/fJWVNIXONIjqrJv/xeRuPPth1X4dLGvrOB5KvyOVjY3RmTmE0s61iw6Q8HGfJ40sC2/jTfR
ZMQ9lRFPDmFFYn1DLZJgBkqQJJnz7J4LXBWgVZKJ/LArpaVMa3WunT5/t2+Oxxzc+eLyv3aV21tY
/stabLpx/+8SaVrQs4OnjST0oY7raeFJ93v7/74TM5BbFS+HQrjpPpmRVrsiCiwWda6OLUoXcVWa
dU3vurQ0Q4yyo0WK9meSp2pz60c4McZDRatJHiHe1scCxa0iQlEh5GG68Bd6TDtnea+o3ZBI1WG7
4xndSg/VsU6qANkw8fCb5SFz68Yopw3+bILRVFCVSMPoWzkmBEiDhljCBurYAXb9OmJoijmBEs+9
ZgPjow8fvF4dufWjzCuRI73B4eyrC8tUlroxaXZwjBqgFyYK6AbTegHWz0Gk9jwc4BW4EQFnJndX
+5jgnwVGIUJZTdfxb/vro3niocw/TGo18UGdeV0+n+pXgPE7WcuTuqtoTB01n7P60NuBvgaxLCkK
7Xro+G9NcyxSa5yfyZ++NMVA4nRm6MrKYYU/pGDGqUP2ylxAfESOQEjCc+Bw8p2Eq6ru1zVYKSbR
KHKo/p+QIiaUcuErZs/UfXvSjohYxj1Hv0dg0pvDgJXizqzhi6RgSl7BB31n4Rps+RTh3gxzgOaN
UPDBG/ZgYfOVZLYV2UYKwNzm2nU+9u+J2K7+gIZ3P7byfeKBSA0JdoQIo7nbPWMrVnmV7K5wUcYx
AlCugJ7V8PGXH4pghX8OlRtTXlF9tAqpuyy4SsdDER0GXnPkiWknxgLBz0NH/8EUHwZeuKOBrxoM
EmbHxCOvwlMNqQO4YKXL1AcXF5ALO/Fw8E4dReAjmvEmZA50rjzwN44kFEQWmV5BKeM2y4PTi4pJ
mKQi/odC+h1U/o6UWrp4NkZfz7p/2IbSmThpdLIH8sPyJP3Fx+X3mOs2MwKoiR5EBvNfKSrLGWtI
PGH5kGe6D9guLTnuZyjI2PfDWFB1bFa66wDbl52X90+Xivop/SsOvED8zIl0zVxKwu8r1anVPyQK
k1Y59/sNMy4OR3LZUqD23G2bAm6NxFYNuM+Z95rqeYGE64cQKqd0NEInuSNG1kyG09kWP2DiAjxh
SaUj09AxMDh4YoHuQ9k89U8JSSiNJE0Sq+2DY2vvc90r7jiDDuH1Cz5ENXj7KTC7fxiU9sTcT6Yn
oYqnnsVGqr9q8gCPRmJ8eqljrnZSfJV+3pv6BG8DgSuRQUqg6QLK+BosTRlJQCKo+rg2tmpBTrhn
pWqhcuMGjN9SrRQIhzrreENk/ThzgpUxDkh3ZQ5/HjmYSDHsXo1NeL3VE4X6beaAFJ28lZ7LZHwS
xDjymVH6Kd2U6bvgtHgdEMvlOquR/AYu179pUVLf/H9GSxq1c0JySHOz22G/UbzA+ZyRgCAhvJT3
WX/n8bu6fzp6YpZcdM8bbDm/f/YwP/3zt1S2u+nfRcg0/FQEujXx9HfipVEIoYY83iUoZRBO+3s+
esDAgRYOtQgXS6uj39cio9X/0YhZwQT0NPxwAZYsKb2NTHtoSxdyZ+U+Tn5mxMRFlmjD1CHqk5DW
dABqZI2mZUFGpCXH08DyJcmG9WMiMlfviIIjVd0bDsUbfurC65UTHa43YNJL5VDwRCIN3IqlOSPJ
75xcZKrwlmtYQVJgMnkHqt4smSwXbieLfEmo3QNVlhCJxE6iZ0JcfoXXOetHgXGwJtM4+Dp9Vn+C
bp3BO3/vSrcc3KTcN8Bqk+gYY+qPmWIrGUF6oHS86OtS0gns3Gz57MJDg44fEPInT5E7pjTe4IVl
5ZXTlxCIgyZsBGNf27IVq8iZmdrefD7xpmY1tTNhIDMjgDTAfYFw4S7lZdfFt/lRgbx71ID7Ki2L
PY/WShP8/0VO/AoEaMdGd5P/VRLI6LUPi8KfKhS2wK3pVs2ElGwn4S4NLZrAQLbb95MyNquomGtG
vffrWIneVLjcklOdGoMdKptqHS8LQOvMcsWWL+E9grGxfNWIA7d8hzvp8lyNMdc4glR9IX1xCZxc
bjP913cjlkwJpscI2gwdsTpv/aROcqsZ4EIVmZmjS9H9Pg04hygjKGgIVeU3U2xk8QOXgqTp63GL
bh3XRQg+29ykjf3tYMhiCe7SSSuylpaxp5mqCV1HkZ2ylWUxuxs9c6OasTFFd0hKfewPLsSIu0UW
QRBraBEqKB6kRgOAgi0edAOgcQtDp7sYvHjxaA5js8iriidHYMzHklpJAt4CslS/41cpKDz1Ol2q
BbMzhwXf48c1eDU1vomf6xFcwUKr9E4t/KTIq5zglK0anFUSJK1YO9TILPmGcm7F239nGnlaoLYu
6JiVe9PV75W04f5hZJnWDsocaBGtdFvPfOf9zrY6EfeHYD2sC/9PHBWotw5aGUohUUaJl8+/sUjy
FENvojpjXHS6O+GMq3ZWQ02xpzu4f4G1QpLYHL2zDrX7aG4UoQTLT0ooBM8wYZm49zw1LKUa2MVD
B38zvNxLpNerNVztn6nHCb/nZyYX2K9KCsiIF7kYKBsz8gZkLqSPvlTUAmLZE5JUBAkAT/F2zXnH
KrNiFxsov3InNVHOUG51Os8I46tT6u4gR96Q2sHWzqNvfG65ZgwvnV1KosW7hEyCEbt1jnUO5EcN
BZY1fgJQuKha/69664m/AP776jTDUR+6M5tIXivI9hvXOBJWTbBwG7FQ+kX83Z7yfHILY1zRzi0Q
uuf3LM/gv7sJmQbSDMpf+d3lyBJ0bNp8bThblfiXuG/CvrB8X57yefLw85nBdJR6suMNoRRfVzoR
47PgV4Mf3f9KwZP02fTpcozzjBZ2vXKz/PqAEz+FWwyl96XmZ+LCjxCm8vnxvePBUswoXmWrChDS
HujwX5U0agdpHrgMNUjkWP2W4V4j0a2pq+9TLEupMzYxETxnh8xNbITo3mKmeERJWbEzhD8jdwgP
pJaw34rVudI80APrv8Dd/PCv/qYuQ+myExnOWDdWrEB+NkblITTHC+DiOH4uHYXbXzNDGv4JjV/h
n2uK/h7eClxTerszkxDoOjakjT5qQI53P0ZWNa1oCReWinp60yin2mzgyIaAm2JGBYve8c51twK7
c9owFa8bX/gu0LmI9ackY582RD/ghJSuo4LEmE6QKcfNPaJd7gl0R4myxlLYO2hGYhxTkiUwNF9u
MnuKHNd1A82Y0eQ4i1awvTPQZ2udrqoixvob/jhUTVvGK0WSgairCavrIGg0PJDwwOK9LwRHNbKk
RUy0Ei23f7Izo5GkvRdl9aJFPsSBBA7SuaauJARbFk/vTaJ/UAF6hXJD6B1ZhWhseJbIoIE3lvkc
RIF5WhXkjYbhSrKqG6zevhnAy1mMkjyOmCTh2x0W8ON7UBAUl+eEH6nXfOOBZpn1K9X1j31GGyX4
+Pk0hAoeh7zebfexAYVufzB4x8DITwwRBsh0qIDXPCUZDkT9HhYf7MBrOu8YVdKvvkugdBak0gis
wNZhGU5ha6gEb7k/rIi1VWp6PTu8qjYMapDZTVcQaMM+HbaOM57oUGZzhIqxFTxlI5Fs5UWdZGU3
WaE+V8uDj2emKAOHFyzvDLybCydZycr13kKsTGz1qAf+lGC4onlyHpu1SlStYz/Q4vMih6yjnaSi
U6uV2rs71+5J6adoZ7A+QRDjl0ds7h1H77DE4KX4hoUJ4APzveDsiLfBzOrXvrBxy70PnHXPU9v5
w0cHeeZdKlsXBG4erjEZohWkJPqBzU1MQ5jmIZKzirwkYyMw5d352iIejyFyt1DHMzQtSZBvpuK1
PA5ooHbgizgbUhniC5cAop2pg6eqBmRavNTlk4Szl3O2Nz4bVF2Qz1Ny7/Zt1d3Rblc48xHW8fNG
fzWcv7g3+ISjuWmSbvtmxqFuHhhbkBsL+yWo9G8/u0NoBgsC6g0zbRP8pJnKwcZ1lqxKpWPVVq9K
3E0oqgDXiA2ZlUJwO1DNQv51CnSIxvzixeC/KPtE2Iqg8NGaBCy0TNR2IBoO5yirKqpz6DgZ/6CV
FwzlYR3zOHeBTPw0SSrd0Kpqou25jNNJAScycYS2xfIYGTE8LG6b808IIQmjdVsMXNPQ6/16RMUu
9/KbNfq2q8SI+tRNOke+j1CjnvY9NS2/Whe8yVqE0ktXs9UfK53B6r/UBC0GEQjrYZh4CEpnqcym
BTc64ve5IGeDwO/YgZnbPtO8yz3ErKBBU+L4Wz4kABDcho+HoYzGZFok9nKZ5pKCuMb4TZ41XH+3
jj77viiH1Y8FCd+fKz/YXK+0sf5eCKTYwcrrU04mF09VSHpMn4ZfToKQgY/a7CtAb6+P1gjKsmCw
pSv45uQ+he/3iKauS6u5w1dFydYfxV42xsEPqviIOzHtENC4BJgE+Fz5AU0jRikiM+skfi4PQXFy
aQo7LGHhnI+I8lL+q8JViOalOTh4vzm9UOp6DqM8e8JCz7CBO/YJiyFGX+tNSTJaDm6vhv02qvba
b49PzWbgAh/EDIXBEp8YUxkF+8VfYO7FkHMWiPccBmoUhQTF28qouFfgg+s+XgbzVuNT/zt9pLhJ
Zt4wy6lrT7fXw7BB1dOtQc3DU1QgWq2eQes62NoFx16DKImnHgU/kSzkojW3hFkppKETYC8YxiEL
kJZhVG6AFUUjOYFPPdEhKXlOYhDqayo+NF5r7NuUdPlX26ojGAQWYmA99no2KI0pmtQvZei/TohE
SPcits+evZM41EV00fsL3gdLB32koqmI7bZrH9DaBHPcAZD62xhlTYpXaaWlXBdx29Lopj09DvYH
ETUqGgDnj5fyD6PxtpAgXC2gxyuknVAC5j6tGVM5Mxins9rEIU7yIUJ+8Do3kCgg/C6qtF/T+Djk
em/k7Snu7CIQ7XmN11NbNZQn9e0qTxZr60AawFqyyHL9d1zkEcEXYMLvOQ79DbRM0YbUhCyCUZCV
/Bxu+0xeWCQ0VzJ8yqXbZDlhwUUT6oHTLVgjN/STMMDVfOUY1sfg2UomfXHvtrFfGcBkfaBHB/DD
h4dacfBgxLBqIepZw9odCZB4sT/8nMdUaAK/LEQDU3GwdGCXw7dpbM5aYGgNNlJeRF+MA+lerMbf
xXuR7DKQSmgSppDqw39cyfl0xy5+oqxq9k2mBWRFPX+aIMNuXdREzmaLrzC/O/2nQYshuQwWo0v8
nxUjSFlAWD7lQChhKp/uZBZ/fNkYEgyb1ZsHg+gYLdRNsyzoBKpZMamCmVa9OMEqnsdb77+ByWD1
G17Pre0Gsx1W6o/28NGecK8hUvzuVPbYmyrzrNm8np341eqAMTNxsnnor1Nl/ktu25vbgzZPYiw+
1+Aiyms07tDh2W9yoH8xODVs01U6HyCQ1ANBrR0x8NtZYVHGmfXmcBEj8XzGvA6nh8ASR7Fk6sXg
yXe3C01LE56l+sta2+PrJKgFVNl9NIhA8EcKtXBizqIwTBPO53v1gIpsGPzm0RThkAmpXJTxu6ta
rpPyN5nuyz5UCSoMK1GKP5ucVR+EXKSTweaNq73KgE82yBYtA6pzfDijDiz+PM7M3FCH4AAFYRpf
lnU5lmQu8eMQqqU7QcfoxG6mf0ytCs6zmh4aD9PiF2wdnOnCxIylh9GfLIofBKwEVv9RqJDvdPjX
HacpautIVte6O53fSc+5I8T3yZv6yGEVS5HR8hrVPNVQpBx78RJXeMSJCPt9luVlmp1QXuIVcUXr
rY588KHWcLzuCRYiVJRligOR6blYBnfO23cup8XnjfIBe2/KPfNuJKb51bLAL5PbgAQcMTi5LyB1
BKL16Zd8VobCiwGP5nVkixdhQkXOZHdfc+tqdjxlYDXcAcVRReG5DjedcEGnMKYSnfsQ3lF1Wvh9
9/fNC6u6v6MihkxAcHpSZk57oEIknWLsq83F95JfeuKmG3J56FH5TcNRY6xa4ep8vVXwoejdHfWS
FniZhOEC/CDooKzlRCJydaVEBrVc0dieKhNrB/J5pNJY4gJ69ZBpdwUrGOPwZ4O4VhLFr8cjYjCg
ODRR62M9+Cb1FxOnqBi8ZNq6DzwE+qYjIPghBcrLnQ+s12+UXVOibgHwISmx+L7XvFU+BnOpIkI+
X/LG+Cpo5tcIZJk1ssXMbluFds2Z/9TVeaaOBaDNsBqD9YRWPlv7B3OaxuBvRjg3laFXPEDnspip
4+/G25b462W7yk5kZNWuFD+YsWpuLEpWDagv79wx82hyvQZtIoG70k/XcALSBMFhwR8O27tKQ9vQ
rLdmccY8pmYWAzMjm5t54sLRg7ZMZlGLx9Aqii8vOmkoNn/h/IBKWCsNHtqrvYVks4LqOng4BAKC
ChtKI9HLYVrfxokSDzlpwnF4N5Ia47OYmPHGbqTvBr06YfMcKidOistNQNxix3Nste0oh4dYFgpr
7zgw6JedsBfRS1qipji1SOxMkN5uQVRC1jyAu4g/3z6PRlZuI+mYxF+bqp9gZ513MIv1bTaPWr42
Bg7HJPwAqSbU0QkJFzgtxJkWPbhyPp/Ludnf7TUgz2VBsf+3k9eIatW1pnQD5XdVQNZJV8gs+ccV
RYNXM9bbUNnmbY3Bj7fcC4fNmW4q7uRlkRiozNYTPUZSywZY1OJC/IU29HC6mXlW0GVJ4q38oWIu
E1R9XwT4ngO7Mg59fg3AdcJWAMmgIZLoG3ZMoKhaLYBqulDxkFi1Ke0wVnpvIv0IuKwqaz797vq0
qm0UWJ+ToxYonPZe75jWNPXMmh8Rlj73+7xce7Y0qgKUwCzsrQkr2iKzHJacH+iAZ/B8qlOxhMew
tK2fQIoKMbRffamRVHbu7mweDk6lG3V3Slq2DrwC2iJArkHXAPm9FKrt5Ql2VQdgQhqXgmZP1SKq
O2Z+CNcJRHblPPACNpLOS0TPC1zza6U2KdCce8ZUTiQeH2nWeLTBEBa3B6WLHDjw6okapeDv14yQ
IJYKALkQVwWwns4K4Y4LVJQ2WM/HUP9NGqzRo4E2y9ak7tHT3zgr39qD3vCydGLpwzE82lnC5fYb
K5wTF/G0y1mg3MRmCzFHBJCRISBLUiejbnmK3Q3F0V54OfsFVsbn34384Nc+bwHizSj8mfhC5dpU
FfLXT8i3AHtsP78ed05rwimbWvcSyrhik354e7YbDFm96ELtymyUfqTFZFffI5JxOv7xYAh9aDB8
zjMFCSGeJ2osj+gsMCo24nW3fLY1t202f/D5+C7+7qH8eXg18L/ieZ0YrHstVr50j1lSgdKuK84V
ZRL7ojpp8NqCvN603IvzEH3htyiz8ERmiP+EzamydQ9OYYzGC8IP93u8l0qPdy+Z7t0XuZCCe5D/
szx8mxNEaGILvl0X/F92HNe0bJJjuNi2MjEvGjj6XjYHc7ngJYeNw/KzoVVgpfb1cfy0f0Fh3gOI
Tm49f10Qrb/ryFzQILFvAq0PfI+C1koqy1/dDlud5gJ9Bzy6HjAHo/RdZPsTZ+mBN0d+AVu+uZCJ
awwhYwWY4pYLdg0xuByKJdVqQx9S5dH3686aCmRcp7S4Jm/Tr8OsL+w8cBSSoDdxaTwu93HyuJQD
hLDoknRsrbum+yPh2qUvuh+8Nney6b9Dsx5IQ3a18Z0Bw3GT+b7x1PocRGFqjgbccTPkha5v5PiG
/zybSBut15ZkJNpwf3rFA1C5eGG6n31E7TUkMnRNypYJuqEI83XZs7q/vpfpG8bXhz7WOHjT1D/f
z4tClK3BBpF0zfuUXoNy6HUyhCA/dsJBJRUCpMB13RZ+yQEywnGTx+M9sfWyyZ1zzPJnXCbcKj5e
sJm9VYFuNsmRHAmI9DX4AHX/Rwv2bsiBlighbiQFJEIwxR0UqTU0JnjG2kiTdxjlGDFrOIyj/dos
dYuqGMWtwsbEZALg438i5LOugjdrhfCmjg4GOzWaWp+7h5jdVTC/PwvHwKfPAdVVbyOnCwGvvP7r
zHd1x+E8QmJj2FMJoiznwhVnN2UGv0QsSv2WBEhU7Nb0t1WMmmttgrnilqFRAsqcHLjaHx8LsXPE
2/Y+JcDAFRX4U2yJT9hgfMXfKQmCQqSigC28n3YcuPRYXA1C7cW3OPvx46I+1aWoz8U/p1Qr0pym
DBQK9ZPFxdL3fkoOLpHX5WRyKXRUq0EJeGu+OT3/kOJ1vcXRVuxn8zo35ivAJnLBDsuCHInLbbgm
3D6AsgncyWFIPARj0Iq6VbVZEtBzpQz+AAsPAudVJWgu1xyOWGGsGUjavXky4XJglEfkpxxM+yVX
gi2jnMvYUEdOsEqcMHySsHpa2Izoa93+93oeTk9zNOiq2bvTStfQo+bqbirO/1mLaLJE8K5ArveG
gapEXwtvkCbtDWdsx2nMdkqvApjejYj4yXQG8np38gMt10iNrPETEXvzTC3TQQRgC9tuMLV1bPsM
dWDcyRuK6Wi60pPkQZRSELpCXIdBol0Iyt5iNEe0furZZPBrxjo1oSDa31/P0/eu9cobY7hSrY6X
i8WP2UOAconGnscqfFCjvkfJt7GmW0uxMrO4tDoMbO8C5tQaocLdksEFVNYJfCJ9k0hdRbh+zy2a
sQyn+dIUhdiTPjLQO9/trHqP+dbtu/5Vq6CbfNK5tEjMpq/Mb8t19awFsshGnVuIc7HLwz8nK6Dr
y5sv1Lp/6lHbahLiiW6fGrRHZz7oursa+rRnlqVhNOhPLwE8nWAtXcl/YXqB1MLbWXRfESMUN0W8
zSB3K/azvpYXAn4DAcSHtVqJaOcFNo6wn2PyML0zBschL0GljifEsj6FtXrGEs/tDqpyg23jh/oS
YZa0ePquU/AmPHgUaAKwAM4zMqIbLc/fNUEO3AJ6IVpBgOSvkACjGm8JjQ93Zvxf2UWrKtt7BEy+
zgSlSCYqbicwfkAVqQNHK2GV54d2803LVaJyGnVbkYn/TyJWFuntovO/DGyiFiHRlFBBa16yqKRa
FxeZQIyWHmCfHo0xkMOS6Y3l5YovLabKxEr53SC6r4a55l7ls25DRNe0j104kp0rgSRf9tFjE+wz
r/P1AHbI7vGnAI6MfK8sGp/KEzIIs9xkv3Jilc9IBQc+Ptnen5O4JPn1WZtQVDxHNYpf269ggVa2
UJxm9pqD8/DLgxAGYVwRXBaDB6J+hzkI+39pasZrA/+k9X8Wldtcf3YX8Jjo1w1xfKMHOet93/K7
05jn8h7R76sBf98E//5FjYG+ilBj+e5G3GBDODtmdYhtOOVdmz1+FjdO1Nsu6PoGM9dKi4WMDx47
s607mL45oQ7vvSxps5kdq6XqfskeCVGjFLq9mbAgzd9/iNWz5PyTgMWbxrqSx7Pdraq2eimjWRM7
S7sKIRcuJ4YeaI+fd6ucpcPiLUdPfelvHtRbAP8Yc6hZiP9QlIBIKP/hOJ33OOEqqzWWm6OI8ojO
6txKt/7GoriZP5sRwRQ0GUMQTvgE5jTVQ4HDZVioJMk22OaJGyoSIPBJ4JIwFKltHAErPna3NYZk
x2OonHWBFbtlFSUGMlvwpluBbxZRCjcyIDBFLgUEl8reVRIXmzf/OoH7bgDRnhGdlnMpaAG0mPtf
nQMwqflLAVoPP0nJ1NwfSbpyrX70EOZd8tKMs7tP4H8jqHHCPulYOSx4zWfVze7JimZTT8BmhN2Y
kbr04nDtosO6ut1mPszL+if/rujvByN3HrIqMWv0gk+K7fWAxkJy5dgwRHg4BLQJB394dtOAfkTY
9i2wJ66+/JitOVONfN+fBc+XNrSJCkrU9D588ySLUO94X1agTyFDNGKYGE1+iBw/AupPyO5EjAXg
U+4f5CoduW7fShaaEnFSdIZYFEMfIAafdRpGgzxuW0FefTm2eUbxWFK4ervT/rIKVQ33qC71HHA+
CORVFrHDUWaz0Z3EAtdBhvma9poWxH2gjpGpOFutiAhP+g4iQep48+y5oLLhdTWDmzENMAuEr969
Zpl9zRlD0caSFQeeFO+uCE3e6yL7mHFQcW//D1w5jdEtd6fQhQKXbnnFkCWQC3nwfb0CIBohRhzn
mSVf2wVwWlHxRZT3ccj8pwV+Op8Ay0b6sGSFNzKnRTbkAOCmtNqryH/Vbc276MFYSnuKAr/PDN3+
+JUqZRbqsn3CAz7Ag8j33bDkX0YLcJ0R0j/hDC5P0dj8micJJM7O+yRZrljQsrczxc2dZ8OSFp3B
idkVrPTJZXXyHWNnniAoFxqzCPkjcGD1rGxKbNCJra6yDHcOsTLTUyN8pzeQkyRpMxL5b67mkG9H
+pkvEyV0+s1tiQjny4gSomO4IetC7PRAtLi6wSVn9kAnoAZMsP59/Y8v828tnCCwSHjhDqhPnyVs
yCrguwOyF/7oNl1SPF/P2jwORmS+lIh9uS92N86JrvxkWWiph+EBYOoSRpsHUrdpVdnbq9bSeb5Y
dL53MgOmVwjXXD9Ky9JWnH2covNwyKzlDJ0dN0Hlv3YiZAzLv6I1lK3LriuCCzW+M22lo0YF8Vgc
I0F1RTZZ7ExXK6AqLCR++b2a/0oKuLKpfcMwXXhUOdMj8i3j5NBA4A0leVrXkg7v6GRcMZDyys0f
gLdmP6D/Fqmb6VXZLJMIxhLHUNcvYdORuxGIy6LrRV37NnALcUW/remqnCHvM5U2Sj4LOqERK2T6
dxGhvdfXpA7S3CeIjzvtmychRbjPeau1SgLJpPaVtzkEcJJ43qEb+ihUv4gmGpCj3c8BCn7l2UVM
8ZB8yrOu2DGeS3LNnPbGOInDeSpL/ycTTau6gW8LY+C9e6g/HVsx+xzsf5u8nkYQnNQpAYf9WygY
DDNGZD2KLWKfTK1/3g7pHWCGUI4y1l46cd93HeN+Esn+7J3gxA9f3p1YqxZksRALhV4cXyR6v7rc
I30Yo0NRtaLQPTDRvTTLeMZf8EbYDirBMuNYEnw3UNiC12TDccNs04738AVXI4NKz8Pjw3Cbari9
zDkbnMds2YjBa7T2gJI0xghW4GP+wkKBK4YreKq7mihNq78ddMgI6UEpkFwhSO7CjXQqyQ2tfIRS
danJwabyap39xJFWUJoVuLprzmvvgh2qcfiVuTgBDeoBHuH/caiznFsjbDA+fraGl/vc6yfnY3QG
UxyqnXqBYE1QYTtcJPrFM4p4iPJ1KMQLedHsJGEP4e9gxCn72tBHXTW4bXs4OnIMVy+4EyOT8F/J
VtfUfIBzjeo5HdZIWOCbVw3t6/+4k0j5JjF4W8Bq87yMTZQyiFpSkOHPa0BxAx7XwDZhQd2nP2jP
DkRO3RG5ESx9edNsurFOgc+pHIa3sUI4mmrDD16msRG8efpRTxWe/hHjeRP6MF84piEZ71TN8X76
40xQaYGMQvP1Wh6/mU5sv5O1PaxzYJZPVgXcnfn1LSZE5yA7bIuqGhchdakMJE5qjCzw74IqU0jn
ifnD6gJG/XgmpAnDeVH5DN/psifV6swnsZtjJ84LVUst7oTld/wzMFH9Z/ft2oJ13qXNfi8tRGS0
zX4GUI0wfi0xfV7VA/F93M7WeexfE/Sg/nhgUKr3LyPsUiah9jAbLIO3XhOwjQN23nyOLMZAGqSh
JNEY+13bvLKSGwPVbS0D0ZcQR+bN5MJxnmfCzlwE8LCHm6kmUhDSdNMLaQHmcryJcEVdIQMGQW/B
pbQXLGS/Lk50nza/Qpz1PN81pWsUPo5iWc5Fxy/ZTHA9Svj6IOdFFNoperEthqtbcD31uszS2Isv
DPBJdCtpDNqkTA0VIWMz5tkH7vrGxw86XagaGz6PGZpDyQmOKOM7uFxXrGKF1H3Xc2aI48BBez3d
6ZRshz3G7gq8ceIcmnI7Y4btY/AHykwYsSqowZF469SzmseW9KaleGl7RkXQhaSSQPvl9Ahstdc6
VMc1y6Z/2wsmlew2Sdxx5gXTPwvnWnLdJ0NdEHGnaLin+FZyjmJb0L7/XoH2DvpkMxs9o4LT1MLP
uH2fAC1taG/Knqw22ClVBdhSOk/9bm8Nh9et854XQwP5rSde8I/e/vgJiGakJOwc2rGrKFW3Txi7
AeRsIhNll80C4mjL8SXEzExlr4InaDX6OT5Kh41uN839fJykhvN9TacvSMsh75nGJPpVRONsskLZ
2wqBUgp4DiLgJw2v6vgYrvOjj7G9BvftvpYu2W8S6ztYusfG8yhlu+PGBec3CqxxxxTDvHoHoFrg
q0aw+Zj3Qw56RcRBKI1iNqazTpU6DeolfCu4FaHV93pB91rlWRWfrNJNs8ZugX+qJ4q8WRmwqhW1
DjAOfz/+m4usKZJ8bWqDXlKDUL52cGjRvrgslO1lU1h3k+y+fkEU/XS5n78+6Y0V3AIEuSMgLkLU
gUz42N7QI29FH466iYKl6uM47q+4Hdw0/6yCRhnPxWdacTj5kWeNkpnIItyKE+cmBsKmAisU6P9H
FCpiffa6Z6eTD3dpDDN7BBEUZwdbmyFT1K/v81Uw77VMgmmg87hdsSMLpbhqFt/BcMO4DdUbTCQ6
BsflRzCn//W/e0MlwAFNMakHQvS2FHUIQ1vQBhNeANp6Kw2oGycL7nZyExeimkHrZnA1YwCwpKxi
JhRYdMv9/dfChq5mQZ1AJBbhPk3qy60Ln+C0PRhvYw2UEblRUki8oH9OkfqFT1IHApnz3mHBNPOv
woXQc1MFY9QB4uCQyyEoUwRO4/OUJY+ZPYK+12ga9VAjYzsPMlCmF2sZ57wkZw7P1jtLDuxASFhR
QC372edqh6+eqf6Zt9ppM0raxyoTQSCTfgFMs2r3KiUKX1qvhwxMt3ExT4abCLT63LBaZR2hlTF+
Ul9IuUMVTi7O85yT2fC37O3qxTr1t1ITPJJgvcv0dseYmsEt/JgJxusprjb6I5eelYNNFT2M5Dul
3/45PhmIzj42ERX4c9qatRDVd4WiZvV54DhvJOAv2W8VUZxp6TXu8+iZC/L94x19cp0Mc+QTC51Z
x5J02hin2JDHWgjYfSUYAdvBStL96fflj9zhQGtMdt30pKbMO5sW+oAubnQT0/PCUQEfZbRpIs+3
BnF9ytzuyW+3HNDHZ59Z/f62u8H39FYCjbsCMsrPnXuW0p6cblMnMengTpt56c28vg+PFF9iHCoM
0rBfm36RTiMW/WkinpuqT4d2ZZGrkYkbefjr3GN2EeSsay5VkK46OrD405ONe2SFVqYq/xRM/ipg
RzjqaKfT5vDy8GCBex1rfSnSDnSU5eIwrLjQf9UxLASgbrvc19neeZb62ruOTr228y+odpDStHdZ
IQxO0BgIDeh3O6XMO9IAamWJ3X8Oqt4J+Mi9eirJiXiOwsQqcTTURvnP9ZgUkOb1twdrSQNY0ZN1
cEIEwO+bFWL7Lj+KYgA0Fc5p4PW+gpi/LXg24TITsmG0nzA24Cr/7zQmohMVebgUWnbTBTQAR3eA
kq+9dfghqjlSmo+KPaDK3ivo9/t2hDAWT/c5LgGAFWL5/+Kv+ngXOAZ7gOhdQBEYjgkgKeGFSnk0
XwHciK++g8E9KqH7+uDRGylLVLZu7s80ga2fgjXCQRwtHNVty7BMVMHyaQu6FrLBZCc8xzXau/SA
2vzd/aHBMty/B562FRT1GcS5HkZc45GF6y7Ed8InpZr3myuN3JwpCCaD2nXgsbSLFG/egPmPq85B
vJSoZ1lYBN1W1O+S50GaHLt84nlZU4+qbDHkF71i1zwm2Jp67VAu3g4ivOcdLBH/i7e0zSitY6ug
+ygPmVzsCPkwZbcmazu2B22w0BWnFpIVipwqoUmBwbz38G9lCKhmggoy4pm1Imtu7rjyc+Cs/dR1
HC4+84NKPq15Ko2lEzWijF/IE9SUJ5QllFFLefc5Zax45o4xTr3c0l2cWr1e73vOsaLuucl1pkVM
9QbDBoRSBvRc8YXzgaoLPa2bF4R4s4KAxDtj7bTOS9MlWNtANKI8luEDvG0p0dxXIuviyPwSYo8C
urmJvdXJHAlB0W9G/APsuvd1KRDMXjtGWUh6i7KrgZr9O5VAzSn5DRp19i9j6rXeqGw1el8ASSng
gv4/AIg9zWPOhdhh+9dEsHbwNiCJye0Pyi49u3sQOZxgrMU+wub7F5FuymtNiLEkaAHTmRwSzcWd
CDlk0h2flJVA6dk8K27gWuv18cRkkg54dilC3CpskieVPrtAExvawJSRzMamhZUXWHNAlusGr7xQ
dfqON0BnsHXz+CGZTfa4MQ+7UN+GbO1yhlWsAl7ytCAZVe4UwNw6oivFYebkf81bnsjClpuxQXuW
KkYlbSiqYUKcvNhnkxtVmjlpN0kNIyiFAwsTRHyyFry7ARcJQx2Sr5DbpxHg1sLs1iFyV5JHB71d
MNBHX5qGfx1w5OAe7tojHSEPHDAqZhobRPriZb0oIsyMBC9/SWwUha3s9DiaIRzG5JSXE2EFqBLL
i/q9WaXn1R//S1N7cdLH5B57twZhG34cPjOAqG6Rkz8pwQ6eldpKxiLgz9kkC3XDGowkPmjbTxkI
ZeAfj05JCZy+LodhpuUbUaGAxaCppmGSWjMc02pw6Q9in27uSFy0vKYrYPVWtqOWB0uLAuWrwv/i
PXTWJH3inNDWt/rBpwEUiqQc0A5tllun9BH9e/Fu9qWD4wHj0IbLQPd1S4J45En1W04eaM533QvT
Wy3WWSjF4LyiVWpluYtccUsRYZ6rFIw+xHUpnF9Wokta8uUBA69X3iGR2OPXyDUeUG/y/RDmr4lO
yshUJ6pnaVLo3pfRsHgGEUSBSAxnMv2w1XgxT/DHt7QYAgyvK+2K544RJPXDKMfLBXxlcZ4CYoru
hnkHUV1jy1WAFE5gDnOoWmbZFEgVI1oQfexuOjr0QFaXmZFkUT+64O/YBcjxNl0P+BLJP8TEmjkI
uDCmvGmZDW16Q0oXI/kSGBOBLaDk0aN4vPThYrY99Z5oIcI0+fcxxH6KYKLzs1unjs29JPcD84YV
xX9neXr+2wdr8avjCe9BAzALd+LnldWPTOsN85D1xMrwf6s4/mITI+yk70kQ5SxHr+BUiN29+1Tb
XDNUtxh10c9CdFf0gGSjhkzSYLa2sh1m2eYksdUw4ndpHIxhP8Uw6YeqJtZQaYAQ5AIjRskkyimK
7kA3Rbj9x3X8e54ihxCqPecLdS0yp49NMJ7lF772+Tk+tqRSRPY2ZhasivNeZNWna/7MiNy/vF/V
gbkWid1VLx6aGEkl3oUQL41KEQbD7HZ4UVbBQaezNsAXAi1YznsKEiO1YN5QXmGGdV+MywZjFP/A
U/xsAxwx4o+5srTHpb9RtOSAjy2GzgdYleZLmmplT7mSG1OMygLHKaJyjoAuNyyZupRSkr+LgCxR
mMQO+Mkj0kmBqW6dtWjNdb+NMIObwALaZ+lMlI9bcEt4pSKhaLqiVHp78AgYfUDXS5laRsTx591g
aUoQUCGBhdwQTckcYzr4zv8rCBmJ6iXI/3+44ngVQL/JB/WuUqabaCp8j6A539U27ZGPLJZf3lSh
MuJo/lT0+9MPDlk92ChwNflE/B1pCmYf1L2IGsbVlznjUOVJMmdtZ0LYdpxRT0muj2A6C4axGkt1
VaqXjgOt8D7c+uONJAqQzDkh2X4y/bwnXpTKYH3xfkiUEoOdvrGlBV6m+FgrmoW59Xc6FLtsk3Vw
KlB6fTeB5fKk3HUoIujr/NUYiOPuqWaaOKpU/T4cX9L0bqDK3ojSU0SYfE/wuNeSPMXMhvopkGq2
5R4nMOgsmV7w/2o0d8YmAa3K9L5wONuCipk62w7dxWVpD/AJhR08GCS82L1vOH3g8ReUTmp52Njq
btglObCg8ouUZ7Vi7uXTT0PZiyU0OfA+qZzkImt+GHpBpuGVHh8e93+Okmts4/nKcuQEUYcPKA6w
3wpMwGrQdNJ5AnQQRGwninOMC/fW/oVwP3kOf7+LGOihoSmS8oclfYjaSk2uRV0AI5HLyeZrjEqQ
0I37qkqMtFu38hUGELNB9UyPHnRZdLgyP4fC5arAeNdKuGX0LcZto/jUAo5SaEFa9x0UKCDLoDPD
laFq5+iKor9QcNaCo7lfiQbcXXpS3ffPqWVG4qF8Anssg6AkZkMeVlQLqRNQ9KhAJDVkVy2mJP0m
JmvSKAaI5QLYPjrkpZJgnbgsdva48Mg36jByjekYLe5gfPajGfT6XKwB1DFf6hiHj+mWqsSNzlnw
6Pbk6mrudxuSde73EM4252Nf2A+JGAJhVapSNVDXzFV3eDkt87UeaYd/2oTuJjfluYQfVU6Orv84
8MRIA0NHxyfEv6TmSquzWkxeIATzK+IAATh41/BwT6ZlWIE81vfR9fNLeh7Fn9XVkyxWAGOUdkSC
axWEwyrvXfGNJQgoiWK9mPvmmaaOBDJml3b+nzfyACshqmgFvLrsjcK90tpnki+hy4AelP92mnAU
uknuJOucShacGssm/sSHoh9EuY/7VAQtVpRyEWCoe8apzxwoiCl5RdoDgRlnKUUdhKsnP4YaIig3
8kwuCADJ5pff8l+iPio4QIFetJSKPsDVN8Et/tCzPwfn7gtKEeoa/1p966Mp6UDqyNmbGvD+9DOK
tP8CygOUx/G6/tDXRZwe0sBofqdYRM/4Ff1LB60rKvfvg8ADVGeIGOHVAqiaTExDHN7ozT8mvAgD
8jpAwTNe7apodZKEAt95Yomd7bOXY3K90A9WLzrQaJzzpzbzKPyztQujRqPsIj8IFz9lH7wPofAy
ztSquihOWaEyQ+mKA25Gz2sEQOvtINphgwHubnOAvdUzZJfuZnAsSKx/b9XHod+VKSIMz4Qb/03G
YKdsBBr1upfF8gYcF1k/IxDeGCpWMzUaOhOGx7fusHBoiinm1qqoM4mGFZRNQ3ynkLx148LRDbf7
6S+wbv9N5YakdR6v6kvzQikQZTb3PenfBs0dBmeb2MdVxINowelCvcji1Y+2sLN3IoukM5lGpvqP
oka5k/mEpHcDZ0WXSDFWFVDg5gEtIEDv0I79eOZ3d2bj4X0+xy+fX0LpNonVSDOstNggsEipS/OS
cJIC7fYiHBbJLTyZkUq7+AuaXQ896l4LY/s4skzEpflCH1F+uyolbt0JSI+yIpfZ1+Zw6vNYFnaC
xuFIRJYvIoxS6r7Jyt+PGLie9UfFYXDOi3KzBFE00smYEWN8zEk/IanGNfGNJMIBBp39mHT0Hojf
C9v56lZo3fp4y//9fHj1hKsL5Hze59B6KU2lQyWLiqTlinpRK0IQGhmKtHaUYVygp5ej7oLuMHNr
I7GygSF7eMQvzGpmLe/HI+6ggU0Dnvn4T+BIXd03Om0rhk41bwkkCtplatIRuHwkkeAZ+4lbOUy8
nq7GeLeXk4oa/CjPYhs/US6CTL/Gc34DFs+/2GpJikY84PN8sbPzjPs2bUtTwDCQBOody52uUy03
Fml26x0Elct+qoVRiQn34YvXiZqNJp01z4bzagor6Sz+XEPKlSHHcZU0Hl5l0hpdsUAPjhsvf6fd
MB1qf8EiPhPdKaGVT8rlc/mvnGdhgFzUSM5j7V/kO61PnpGen5GE6efGgUWfmLRa55pgY1NJnrVo
0UWOqumzd+wiGyBjr2XJboyxpXLO4JjpsA/TN3UQTJy3++B1PWmH3RWELayCkQn7lrUdm4hD6j3+
4g4EzjjYt++9gDOmzWxfSsNw/85s5Ayca7a3R2ffBH0QRg9EQ9WsRAqtDfALpLVzLRkruhYPYJcB
K6SevQYqKlFlu65ClTy0yuI+TX+z5vsNn/aFou21MMrGXW7hBJ6g3/1MRYcEUQGC7E4GMwKC9DWm
HxJ0ve9SU7ZEm7DvNM8a4v5IyraYMXmlioDu1yuVzPjV22JLMAWIR7ZLiorzj1CTDtX3tKkBdtfI
eLlZ3P+wTolJYkmKm7N6BywE7SLTaVSfZ+5ZL9VQlLr9pXJm6ljtnSxh8Wha0SQuYVj6mKwtVbg+
B7lA/yZ8GQhXxEsvgtFp6OykjVBfGOwXGjbCkhSmS4ao7xOzHjSC0EFKyFiyLCPBK0YqbD9X9+Qj
owKcNMhNcn26hbEYvvWeu6v4FTVpm8QyudF+5T4m4XlmHLyLxhSFyKvnW8hGL4E1U5lkb4x/EZ+d
7iDk3mJwXeBriyfErsj7fT1NX4Xd/wJ+X443qOYbaH4tJMKp7uXZTTFOMATi2TZ92X1la7eLhPi1
xTqiXNU0cFoe0R+o73Buinv9TzOQsnEOjaNHgPg5BZd3MmEGBaHFYYtt4mmwIpbaUKrBthG/Wydy
If6nFnGXZShqRb1/PJ2DQW1F/bWyzxQA2GEt6PUcxKDVEE3lfoSATxtruLAVUX2zxZi54r3JkknP
pOoE5GfAOqhLST34Q3Q4Qgi+lM46upJpb3kdVEroxHXTn3MLGbOUsLrLix5TOJ/vJwR66mYtp/ll
C5bCwrQ30sNbS6lsjKxfnk7ZhMtGiAWuAkjqiE9Mtp6bB2+zi+KFD19hKqHFXUKXHfL5tnNS5riS
ZC+EIt6jPxmP0kOoySZ9u8fJ7+CCsZk2wCTlbUkiAbbmTpCIqARM8Q/ULOhHB4hXPornbJy5dbFv
N4EZLl5knBCa/TRkYICX2A+V0P3YDr1sAUnrbLzrCLsAOQ/ogWoUcSrWjls/ywI+Ci6pdowrDqmM
JU0m+Fk4Ddq7nc8L9PFYdIH4/kd2KAOy9fNQx9v4H5JUs5vNytY2hQZPzbyVJedyoteZDaL/+a5L
Fg269PAqMDtWr6Yc6/ZJRKGtmZg8aFlOclHlsyTNRATT47O6CjAbvX+Q+I3mwmszwKzxEhpuj3Ws
HqkCciTMV3CtzAZt19KdryucwGTHMcJ0JU+Q3Mt5u5N4bN/9UnG3i/vBJzJ64z9a5U+chb6P060l
d5JePxMW6wVsxakjz74qNV3TVUIzdSvgK7jDsQaToJxF9mqQ+pItTdN9fpvAOgh6y77b4SMr6GqS
GSqaHscN7a59NC/dTNTXTPnUlL7WItl4aOUzPWMPjzSGnrwVGfgzTqFqBQgsc9cCJ3yo44LnBUwf
Jlr083jDxWpOaxqbfibDc5a650E2NFOUXBDmwD05/uzFpUWs+pksm3iU2fMuxAiontAQ3MIK3WB1
o6EwPo9Kr0YWoRrfkCDWg7ZkJhUi96azMWElaVRz04ssXh4TMKjAoT+L5rTWxah/xbtvWJNFnYRh
IsBLAECLa4Mv/sc/JH723EOc0js0WBjMeetIrrAG1BRHWBvbN1UN9YcH1NrViT0k+gGSFTOwkL0m
XbSH+9Oyg4IKXPyNVsqtL+XxiKeCw9gkFjk9NLegbas/CrylKMu++hTNwZRw52vhOmFYd/KWBkq5
b5vzpkh2PJhVrqRaxSneO9VLL03uRYs5gZglG3FSxj/7CXSihSWWDrt8rO6jNOnzVZZlLfnOO7KB
NcviYhjYAB+Yi5aENwwPU/KiVbanGuAHaVdeWIp5jhFR5jUzX/8F85nkCaU7nBlbqtTjedw8fMdl
qN7N34hs9ieXVuoth3JqKCRiyGYvNlauaDMcn38JvYAScdKVe+XnSt6rg1mVZLQDePNXdu/FNecU
tCal5ybRC2PJjclVBqePPErkOjXNhJvVqgz2QBiHq2BFBex5K+6a3P7r3zSOcJiHXAeqqCkxiHGC
BBVyBWw81CFSn1wHr17zGR2BY3wI+9ibmvHHS7nocfUHan30GW5+z3K4AL1ZOlMoSjbV9faqogd6
oCuqCDgWlWTNdxrf9gFVPjYpx158EDP5+gZ7nFEzX7PPJeqHjX/wWYN4WZqRlrSXcJarr1pbqXco
J1gNRE7qsZrknn4CVnbvfK162UBLhFdIUAhfP5dj7vXpCzQ4KcmjgSBtNGFAUBHsAep1D0wRFmA5
fjNvgGgsd1DBNwDR1DAR0/1g65GAeF7gLpi68jixk/zds9DtHBSxYI4n9BBgKSI75gv4i9M6n+fR
EqY7XXJr4Ae8qLpN8LfTlGVmzbqKj1nyok7k7/JWS1T0oDAP+sYs0kuTwxA9khs1IAfyQJnfQIcG
qzKyytP0Qhn9IhDfWn1wjpo+kRWo4UZFZGolx+UsbOW3gTR0OgrYLtA5zX4A9acTcx2X0ShLHjHS
RdFU52R6G5muZE1k8696C/X38EEM8mv9cR0oOqXNMBDWO2pdx25YpzX0c/kMFoIPPgDItMsYgHPx
Zlplx+8yPDUDcasYKwcIlNjI47fOciOT0G+vtlptAAIfjt+w2yA1zTxzHLKiNfjVPk4YWtUgxIr7
3dtG6uh+cGaOVryxx80D4EcaFl90aEdnbIhaBG6Psb2Y+ID3X6d4YCn+8piH3jM9CsrHMINfemBu
TFrAeHutkVtCC/5FmINWY6wUXtJEsHYCSj7J9V3VpQ4lJW773eeFh/qndR7GaQkfOm2sxI2V16Lb
niHRyaPeNEUee57VO804iTU++AoY/sJ9Pwq2MLcoLrDF9olfobHiWuYRzxF6GdOoaNTZcxVhvEhH
eDm/AtqlZvF5ba52QAM9ffddDpEN0Z+3HvmAeYhwttctwBHBX+RspVmxeVT8orkFI8TeaNV4VceM
LOgtg0kx24sV8Rxn5Orz7ogtbY8psZSHxf8bTP/dBEyqbXxpO5rqO0i7jc2mvFeREyKEbpNJvv2+
5tKSNooBsm56xJ7rhqgTBB2JkFGLfUcGKJmQf/6VOHhh5hBjKOa1VvdE7NIBG1hTVIl0C0Fh4fqR
zVfVvHP+GmtkRA8HKnohrp3/fC3RuumtRgXrLfHoAdW3F80kyJon6vpIoU2IWsZWL9HVpO3t5a3a
PVhk09XyqpYqs5NvZENgJFkU3qkj7tCXzxVnZ1UdOpcaKlaW+3+iL97wJLIdnsKJLW+giderIVJ1
vtlVm5hXU91XdIV2NvKbtowDFEfcIZCbuyrLyuPmfHNRBP9p/r4YSl5GQROZFJ5dq9hiEosERIoj
tJIU8V8tXAzSAe7rLEujjEYCoeQ2DCK50hLGeCepZ1tIx+2tX9mXflQ9retpG/yG7zTv0LTF7iNK
ZKpGy8w/N7rOLYkMOPqGslRWlOYoApqiMPwXNbZj/fFskOKTE+pa6hoLNayIqjjzph9N1CaaXVYW
1iExrkSt0D1haK3HDMJnnV0o00MHGYfI8l/S+Jl5xT0+HtQicInNo5IsxsUsImsajYVoXBxfSs8n
BrH2fGFvhelOF0Pt/un9x5RqZcXbkYRlR5LKw5tCkHaYtfMN/bXV4N/WMn0vhHu4mReYcAAztqOy
2RoiVHtdWRB5iL6Y06U+QrN6wvTXTumGZ27oWBgvX+ua+/NGAxTBF0SygU46LI02gLU6nztV/ZG+
DbjvBE9qacmJa6tgGRX2szpVe9dVZ40r5X5evNbkjNQL/+ZN+DdsJgEO5/OerSag8jkymD1rNx+0
ZnqmDQTm7yaEaZitK/OBTnkx6v8xSFU4HurYIkWgPdAm3CItDe7v6/NUfJV+zfCWYqFfDwvnxWcG
HvNdfIT8XmN5d5xP5kLFxahr+So+CFB2j4Mt7xkfAn2bKO3CpYguVsXp28go3e3GLmeCeRO8mirP
gNrj8oCs9buzMBcIrSsSW0Jf+VcOnhSTma8gJr8L+IhvstRP+C0BrPij4td2NPu22evLlynhr69K
ZzWBwt6vSzMqnBe7TWmIHJ07x1KIcip5T9Ntd8CEG2IGGq2BI4QXxLd7olIyHcGoTgtKgVuv5WKO
fLzxNQvM/RqNWlaiwqKk0myjubysm4GFHTIUp6FyIqFuEIvGtNepFz7bUGECIWzhcgd1q4ZjXhTA
p3Gwhg1SrWLRKNTqTlIBwn3QBZCRXhQ/2GAkWgowvgUICPdRjdistjY7Tg/4HwkO7CP9TTy8gLfS
KAYzFk0HCKHeT/gnOE9r06LbKCsJf2/nn0Y90LTA3/641NmxSLoONy+JIc1paib8Yi5RM4e4oVZz
bF6Qu6MkJVNUY3scaSYYtgUima0KIUqWbfxfiPrNwd64hbL165NoFKx6FXzZt56/MXaMgC2JT+rc
aRPKvZKcOu7o3BkqPAZsqkSXsGVumD1fDnAhL0PekGIH8lQhlJqen7hoPox+OQfoGv7Oq46Qcrkl
jklyGH09n5lEcXUXl8A8D09s1szsZTkGI8e2auF2JaoWqyDLJxY00xyijWxB2JbkIWF7v84gI1Ip
XycLPpTdByMYfcfmJtPHdqwQx+rUbpRk6AU8tTYxz5N5MpJPtqR8AdnmgLCcuSJO7b2y4KIsLiWf
YBrogHevwQMMNCX9SdZowxTie01bYOJpzfjmiCPTRcRhnHV1Enh+nuhgHbsXCCJ/Thv2Fljzwngm
kvYYU9y+GGKehjv9zndmHFp+ocQIasBcpGwbkqvZ9sO4ydVTyo6KRmHCuM4c+wGbplmMpAB/58yy
nmBVUfMI08vUO3deHx5zKvFc8Ku+JRLDYNbuSgzNKpjHpIwSpCdhPO41wwrkYofZbg6fSueUByOk
hjFpWOwALOlgMrP5pXdCx0SxdMNT3v/RFddv+XL7LF2b9/I7PYHQSPWTJGzPYS5lyz1GBdXeSVgQ
u6gBgRR4m0pN90T3SWjvN8cUusmG3YVE/0ar/n2bz50REifQ7h59QO0jIHTYBAqPFmaL9O7n4qxb
8KgEmKliBJ3lDpEVs1+TlxuoG+Ca5vANGDzSKUvmbO3WgHi2lmzrYtZSrB1hr9w8hD+fLb4AVuMZ
po7h7ZeKWIOY5NZkOimOAeOsai/3qL/SLBnFF7Zfc7gREmCYV8PesB+NsldsKhaFTiWPiDWjADWN
kmCsiIteQC84smCt1uDnqBeQ7oN56qLjkLPZ5YiDWKaU/INNpdnl8DmpwI7TpVQz/1dFJHDZTUli
trSLmbX1tgQt++S/ZaVSzf+4qBzflcUL2FrkIvvWMxiuqccy+0RESUoDidimXDK8aBZ69T1T99Gw
qp9NDOELBeIEiciNj9ZgfwM4PyEL72+P6E2uy2FddV93FPSIVE2i6nBEn4eC9TR/Q3GRplSS7Obv
DlAwcq/3e7nAZKNkxONzHLhoSbP90rtYOn7s78FZYGmnILF/8Wbe56s3+L+J1gKDHiPDBhVgVUPR
awf4s2nlmPJ/P2ZeG6sry0+A/PsfmpPrl0FGLlOuQJKzAz7IVg7aVGzUqWM1pe7JOraqojTt8Uhz
hy2s2Qf9ZfyHHSzxXomohkNqvYTmyi9MZ4MIpLcMMPzpaKS+qim83SU5tQcCG94ylfZmAhULCrdy
OvP9ULkJlGrvg3r2foYG4mkpSyP/QN0jO3GPWySwtHWyMV8jhn4EW8lB20EXyGKfRo2rl8LlTdOO
lt5I7DFreL1BfaZf3hGhJBc9QBnTD3vuvqU/pFoEccuPfJ25eRccUwhXEYFfGzSrvmqC7xRlAUBG
y5ruDdibYQ4hhiQ+nDGWgBM+LVIomF6L732NcqjvvX5c+Gcn/BU4/CgW+wxscJ8OJ+B4ZnRHoQ8a
ApOU0bIzBZXno1heUq7CHwGERVC8AbcQkFaCTdYPcsBYIvFsXoEediQG2zF80xb2eollrjN6fw9c
OONuLecajP0BhcaXJcLUV2Hrris7GB03y6vY0I2syyeLFb/Q0pmX1Z1opcFiRtHOnZ7UUiTPmsRr
xUgkKAG9YvXeu3Y2i/WDO8eTtJI72u+xXmqMnQSzNnO5OYP2mkJ0lr1WEz22hzSDwDP55AQ/lBUw
pRCCKfn2l9JrY4vt4hSo8ai/+jYY8fZ+HX2k0qD4FJC1BCOl3+nvE0I2PCYTpiBL20myCUlGEWol
7BU5PTwMaeG9ZRtFnQh25gekcwGcyQZy45T+h+eWBbrSBACVFvG6A1By7Jeh6/A383U3F50sF6wQ
pMU+4mUMX++ppjkfMRnhOlETiDqQWFJOE7YvPcmg3JF4V594+YpYOOw6RcIWGKaG6KjZd9KF5N0T
+jV/5aQNdoYDhGM2YYq7YMQE7zxEka7c1XhTCOqWgrYP440qpO12pRADfedgf3w29U6xIhyc9wIg
eEhdx3j3bVWIASmlEOcFlymqP26UxrgQE5f9nQ4hUj+bvTkUXk4xVvoMmBE1K/ktykYnlafshiAX
5dGd2XZUTbgPcpHwcdRTIVFumtFd3VkSlQmqeON9qQ22n44HLVymCrBz9X1IHUwNJncQYhsPD+bj
1gp9sW5nBKw3e+CBWrlRZbrSDxhNxVvikzQnfiveSc97sBhwcQzkyfKJZAaDmoerVHkdG4PH/1oP
nRa7aFvCGeTOJzX2cv8mQmrqrN+k+yK2UoELatfgiu0SSd7RnE0XiGhj1Xa2kBUEqkoEGQ55CzJL
z2auYCDNHoDQiLd2M8+FPfVyiJKV+gEgoLrCDM3MgwxZST+nSbdbPSWUWktwobzoZEFU2dm/PeQR
/X5GZ0lfcHOQOl8aHmnb70VWNEwCH9KBkc6sau62SBVWS6CoZGnM2DYjN/tNj5Rme4Bza7lI6BM4
mYS+5+VcnEBdiy1JlIWz9p6V9rCEapuJizexgnReGGjER1YZsluk9oej8ens4O8Razp1J+H5fZ5L
KmNnJbFXiBtBmfqP2lmvuJq/U+IFpbKMPp970sD+rAT4McISC0GrGXQXJsIBrrsk3Uj1hfPI2Vw6
/onOdxVrLctlMHuVWaEbMWal7J1pyAg9phrRBlvA4J8Aue16CXV5XNDePAwiVrV0LlG2+NEEZXb6
TxePck5kT6Y20GQhryjIARGimnH+lhC5cWUefwa4hMbw1urPzeZvfvhibDncAiWYRypHB7ENUdYc
V9kpwPUouf6+AKbvad/Na6aHyU/+ueqIfdnDQRMuqaePfro0vVTGEe0KEPiwIlq12FSpVQPrOgjn
b7r9f+ItDOnd1YYKeC8cN2yiyx6qf4Kryd8G0+AnkncEduohRQA1mty/REroP0Yj9ln+8dnWq3zX
m0jXYiJzh6I+n0nHWHSK5LTcCXhZsuU8QQtkFzkyQ1d5FFTFl4BpNk1R3JsqBzstfI7NcEBbP9EI
ULIF1R0pJAMENM62Qn7c1LAydsRwMDwuu50ZuOsVUCzVMC/VmyUQ5dxbVWhwUwjwhlAGWUIO9cQp
AhqushsrJUV2sFVdGhceprFVyNE6PtMxS/QvPrWf3fs0xlS9TBbi3g+B5oPp1MWNwhtL3FAWjkbH
rNLRTzuEphUbE1Ew0jfVBYxm69jrUSA9lpD9/5ZB9Wp5xyy83a3Y0DnRiP68sNXyC1RniCZUbs85
tBqUNIrs5QWiXmVmc2/3rNeCzPIBcslpG1XYkrYULU9E6tMegWgXQfv/gWlTlQt8qdTdvMxayEcM
Gf+0dELUROf2o+P/G71ylPYWJWVS1mqeutDrjpHqvT4UWfMOfaMvFyU6zotyBVDxE1T7T4qgUCoN
WdJPwFB+MTaK4kmr0FDZYNV9f1ViHqaClCbR5FfrNfbkr3ATu3fS2cQqm+/YZWGytMIBNcJkWbsk
L2whOaz+T6DpAjexbYYIa6Z1YH7/nJhf6CNOP51j12E+4Ts7zMZS6+EdIamQZKLbPVESDSHKhd76
U0bKSyteA4sBOGfFAuStwP0W/8vSSxMN/VaMrzJOqz8wqlJHQ8dmSPpF02cS9cjLoTyza0P6IJ16
eNyAoDqPXA0En/rfylUu33phjxWERSIYSQCt8PPz/8/Azcg5LpWRIXesbsfdCsyLlOVuXgvrZ+4h
3/UoJO+cQE/rJjQ/iMzlg4sRrp85VvV5FQ3/aL85aLPnxFZj3UdqzgDf5dRY8745hZYtT2nHwXeM
QMRS/xtAxWCKWJcTw2eP/976WuSWjFVNXRlGhCOl2jOYBWok2Bh73z/5qfQmQDYyVF69CzifqDC5
5VCWRNYZAiJcm9W4oaYjfiimMircw4AWm5pmQGXhNHoiGMW8Jb6irBsEsPKA/K4ZGn9SyX1AZZqa
/5A2v/WBz9dmCXPDhgnRFxylk19scnTz1S/BcIBlzAMM9Mz3tFMQkSU+AykRQ7kYpeXvxJat1VUI
nEYw/RxakM//ZAm5nlRejjLT0EeXi4vQxFbZuICgts9wyJVrHOv/MkRpetNlPXXh1RiEH3UaciJC
DWRL32WLJ5CH8chpV2dnQ3NDj5ImLwFPdbXZjWIGZVV/n9RtK8ejT+E+r2Bz1xA/aaSDiC3F5IyD
srGSvEb7T4wEsyG3w21knbTPJXXxuL59xehAGatgjglMnI+wkbZKyR0m4ODEiBx5qkYYs+ru/ltp
DoT+WKrpiAbaj/I6wZK7u94wOTkW6kNtKUirSWZ9WCRPASTBFiNV6oJZ+4Y0U1KYgZFcOxtTVFgz
pGe12SURiG++Pxib55IJZ/8fh9DCIpyAIFGkML9CQ0uWK4+XCsVdg5KZ1iRE3RhRtgF3hCB0nuV+
+9PdbGabn5Ga9U1PePUcSs1Uq2/gWjcSP0VXOx8bELi1HJpIddhGYbwB61nagvmBW/0mnk7e0cDu
zV1HvmTQIWXjCwWXcs04BkcmVfLjLyiGUCoVosUmaNpOqupFwv0KUn+Uu3hRatRO+6j+xsgxkYwr
tV/pdaFizcZhdJzSyTz1QPcS9IZXbriuErx1IzXhleZkjezejSd1qj63wwWiDeDvTVeR2igC0Ew4
UbABlhR9aEiP+8V8ggkcyQEUyPvZ923SahePl0V3IH9lqFx23kWG6K8m8gLfvlrDxCOqqdXM2i+B
NRNOCrU19Q6oY5O2Gzj6QwGcsb6UywaTAY4hRLOXJl/VQB758GGvtjQmja1hRnEz59Pjy8Mk559I
S2BEBSypUtZ601Vo14zcr3A9+ieashGDEsWOXslVOSydMTCQapeyBQXqW9zyMXGQ0JzaDHa++dCE
wCQnVKeu7qKS3u/AadV5iLbG2UTZxqTpV7ar0/ZaHBReXxAFyLqmkJUH9rxV9pgQXoY7YVij0drV
0BniilX918o4Io5CvnOFcHJozSAehXYkL3aMWxv/pF4NL4dxZiaPRHZ9NS543sbHQ12lpVcLRZ9n
Vxq7vDU9ZN/BQb+nKqXdMOLdlr7GxtUrc17D2Ok51y0qcQUj+RGixwDEmdw6A7Kn0Z+zxeFgBw1y
4BYGxY9BhxAXmplSmvur1+1KrC+IilBRKsEZeYqEpm7Y78Ai48pf0xXuGe2+CIt/y6sYWIJ3WDgd
/QIYmu01nNBHX1I8mBUnWD8acn69HMqDqXsEGF1B4JSVycs6TrUFqhenKZod92d2tQqE7JqcbXOm
n6UDyNsMiOoDH7+eacBhokNTkZSy00B7Vu/2EvYsnrMH97sODojMRZkW/Fd3PN6x6apOz0NDMxwv
hpZRhXFvczv8qmlKXXsSeEJuAuqA1VfnOgDDR+8ukZjwNcsqDHc94X1sSAf9O540ODpTJfTrGv5Q
stI5ypcG+qs0DDrsHTIZBO5R9O1Cvgw/ConkFqFi2knb6D0bzzU26MHPCeAmGfwX0DAsYMSggN30
ZxPSRZ/lWL12WN8zn5z2KffUKLxUyPGWBBrCHuKqDn1WY3lwfaZAY+1WKWiTHqfAaoaAgnzogfc8
pCqpXnq7CVzg8wkxCrol2+PsnWJqgzKtS4fUNIo4DKxZCUG/EZ7aFmqb60dYgGiBjaBLEbrp50OF
8ZGZYu3/Azbm4H9YPE25xm5y5WGntne8VN+R/Gtmuy3s8pLoYn11rWpL5qkSl1EfiAWG/ttUjytx
GiGnoAAVzcmlKvhp1gbjIB+J+ZXddBXKj/06zEyR5s6e4xdFIF8gtm8eQdXyPSyDaink6uo9O/Kk
/UVyN4UqIU2gab8JwGCbpFgTCSbOUTSxRquNNcIxMpPw+pOSKzKkIWzW6kBjbKvR8pco3nK8prdT
FKlnrr64ALNHripv32mbFBMgJnMbVscxOZJG3Fikgb1JxwmhOnzqqO3a4oYT8gb0RveYYqsA8sFd
6bIg4fNIFK5OQSTgtSdDXGxxhKkiWoBTiD2N+Nu6hbTZBsQUUfsWlo7wJm1zKIzhg1qpJxq7yx7F
85Wl7cLYhvRTyUKTKJscOWqGA7tngmWpu0oh5I5sL80g+/Z+r/tLIEq+1t0MMOXX11Svlvm5n8rG
exgp78Z/t8QBCjO8MmbB8OBEFEF5WWfozGyKb+B10EGIJG6ZGJu5a+jWeuZXIFblzMEoszDL30k7
xGaJC2M+dVlgHHuMaso5CxTKfVRDYy+K7FW0XZE727L0E5uRhca2Ch7HNiGIPIbS9qeGo249X27y
kgR/y87KyhHReqRHkh95jRxKfsWtSFwMiX/I+Gg2pi1Vlazu5URIL2S/Bo6/gmXi27dvCIctvmb5
0d/zIadQ754xBvn4R1mJ8gbgGgJ2u37rCPSVxfCNr4ohhwlnRWglVyflDM/0kwA8CID1PMlbXY0h
l/t92hY9g2OJFWjhDIm8HCRi8Hn2z977AMPqF8rG387TRBrzjhoLu73yrUv4XEemsiqyefzWzwqZ
NJxhWMFOaAAnyZvE2WViuxZCUEeHLSqqgXpH3WtaQTTabrIsjQRHPX+Rl/mwILNA3A/RrnLteYzC
FphZw4NZG0PprhExFW8MNgIuKuubGvmeAQRaYqXVpzW6XyJLDhDMpi78GX+mRXKcnKIgLig1RDkB
1M9tZIHukzsbr6eVe6KGMt5oEpaWx3wXn/Ds6bXgw31ySb/UkCBOoYR6O6RgSN1nT8uIUFxptYBs
ZelMBkAzVN362J8Stg+OvNOVtCkVznxkfOoouJeFqgGEWtGNBqrOYedVoOOpb6lIAcnd8ynHIc8O
QmYBaGgN7dLW+lP8QWF8tG0lNuOWPtoKGeOB1jnk2J1XuD6xI4OlvZc7VTiVNroORWZRVQk0B7LJ
LUlFC5ZQ29YjGiRvSrvn3+6QoJynJAQWhPOKMD7/qGh9saXA3EDWom0ar9Nxo+PKZhaha8i2w3TG
S8F92es8yalwELoMRX65ju8eOEKdXu5jzm0AuYbp1IlrA7fCteBBOj2Zq2bfoxlZx7qN/IUp8g1g
xmEojV9+g+5U5YXUVm38E1fwoAwXL+nmGEWHQcdu8iapvtfTgbkQIhYW8CXTbMAR6bTb6Kp1UrS8
cha+Ya/sJMiWqDFGjr1lNPxQeemXPl2MiwW/iNavS5Z7AhjKQVtO45Y5yJDvEmJH1HbfjaWYWBk+
XOzOmaHskWlGFeNYGROvImOrg+Kn1rCLikoy0p0c65uuk9BG/vkwq8+m+GdKw6dxP+5oML+POtmp
fuqF2XBr5Db3MVJeUSeMD9Nfo/e2yHu/61RJ8IszMkT/t7QmNlV4HEg43br/m+oJwCCRMUPLcVZb
hyeva4SpiTY+fjfQHtj6RjK29MNY84v4andf9f3DwkfirZFWzXsfB+ti3mV4yIuwZ8a20f4a3fCm
mWuLa6Iu2HHC/6UvI440gFrQprdhLkjSS4M2bzp776ykVS7RyNs3KrnA68Lx9MYO1MUk82MUSSzA
VMw9zfr8j118FKOlyikBsm/huMMeVhVsH6YKXFlsJbMtujWwTQ7thw+fLN0M+NbLToyEw/IXQceh
7U6TTL5BkOHm1kBWv/+2M8NCL0VUD4MuoRaLp8yVDex8G/kiQItI/eD+eFVSdzUyXPU0WKGXX5Ax
RekQ6ytK+zOeXj8jG6G4hh2ZYSgXbKicGzzVM+erFbfeqKa6SS8oSiI68G14w3QgQnZJxw87P8lB
6KMIct/fyIc5/s2+ptiz1NFmSKNQhZ1b+59IWV4crhbAYVzmI8oFzPOAjZ+wo+PahX5B+cQMY9ou
gsxowrePflHsuRqQCoHW4+eUc5apMDXP0hWLB0asoVBXZ/z63K4U2FcEhcesBfmWViNg2Xr2nEC8
Wrsr1Bo9v5KtExvyt5x/JrYq8MtNJyG1uHVabs9tQWm9KF65HVt9nPgE/j3nh0OhUlvZLKOyIbey
3bEyKYOp6CvkGRT+9DIjFse0LWtCcOf+41uXaRLWp3Xx6ifzeLmUZuN4xveJ5B5dsn6cYmIgSwJS
oKClZnmkPCJoDzZ7rDVdOZBHmkcZ0TsfHG3QkKmICuG0VZnyJu6hQthUgJWkr0+hpE/hNZQkhUVp
f50cEgsnV9lh5TpIcEYfM8qYz0BNnbCeXTN1BTTu4IWWp7Dur/rGvJywwrVbecTVUz/K8GzGFIDI
VcvEi44vnuNOyTaTj1EfBJ3uryotauUbk8KKfgBv2bHhHfu/e5nTJLbZmuZO4b0H0Pk1sw7tm9d6
9BeSaUr+GV+bJZ/KpcqqHBMBqCYEHIExrZev4vcttD77RJJ6HF0oz4Mfa3E+TqDKr/f27r1sfyTf
JgL7Au4hqbj/OXGyWme32LwXWlsfnOZ3FZURzzUwe6Us+UTg0Ut94KCoYlfdpf+EM+j8krBcyCg3
VIXYmjhCuTqx4BnzDI/1VdxvuVTgr6zUqu2+pK2uyI62h2FQDVWCqER8lyJ+S/Q/P7Ur/JmozJw9
vVWpLyhelidGqdtfYJfSBNyHne4gMscVD/5VRQkHV6Bn7fm9Ja7+JB0aWtHzqT7K2FnuT/zkfFwF
S+aJp1bn1bpIcW462JJKTnPi44dGWwiJ7Q/P1InqNNHqUGpDjYq8BSBP1NUdkSqwBk6aDz1n/71T
XQ/vMHLUvfzaRg0zFELd5zUokts87Pi+Zc4gSA2D/Hhn1HG9qtCHtN7e5t9579xGAV0roD0UTY2M
5i5cwMw1sm6XYvsrBB684qLnPGLooLHJCM7/FP8TVX/FFfmhTcIE6y9Jfa+CP3PNbahI1/djsEMq
ptEI/HhqWbBR7lxv6hJ5AQkBBRVss3hpnAL3xDli7MMYB1fPUAfz7cArb15DvGVU4FsfLLemeHN6
7Mfup+U0XCufM0Z54NkWPeehiO5P2NHaEXSvyYBchiPKdOJ1fcTGOSPXV5muIPWOhyyuD8R0Y9DR
YKfvgUIeHUBna2ZQmqxIke2oMNqMnxcf77TCk+EwaUdx34WWxe74fmxGYHoQFNCyt3Q3OtOZcc7H
PFw5PYWBosyncOGNwITFvL2nRvzOGrXSg1Q4Jk9I5zQgCGg/Kj5g4s38BZibCm0+tFzg8zUoVi1l
szGhpgJvFODSSSnc/+y4UBFlcaFkoY0my2TMC6YttGDcyFfUWLV7Ssg0m594oT2QhEB7ydWZ+YGi
BxvZ8BHsQME1HOxXGugj6RHzQBUwtOZGx0s52VlzJdEbJvgNDGCwD/bBpwKhrJ1D3y447qVwgQzE
uhpuHoyv/QzikwSasDh9NrLYdfdoQ4ZwZHdSCimNLsamsKkDGHl5mBs1NWiMF0sdR58hf4Yr+K98
wBdpTkpuzPrWz5P3mU37DXICf0Hfi0OZL9P6Gb+WxtxkxIKrmZ0bFiNm/OJICheIovTIfOcGao2v
mrhknw96aOXPc3pnfDbbCTxmkNHJqFSnl5+chhprL4Q8EGVoQf9/RDdvRXihPWd6AR3Xn3l+lj29
Y3jDCpql+BKWTzctevuYgVA8FdwsWGj+7frDaC3exgFrY1/ojA8Prc5/0UAk1F+x8bP1ten6gnY8
Rg+6uGqGtbMWdwlt9rgiPaMCbZT/jLlpIlBZc+PhNGk1aZqOMqIxd7wzAAQ2/K27sGmV3VRQU8yu
q6TV3HoS9hFca+YpPCXsNEII1L9gas8dRchgDufYSI9SgSMnKNQGoxkrtSDwY+UyNaRTfbAth97x
xsI8JvYjt4jbMNu810mtro3C/Tr3reHFWwAVLu1xc/g1mBxeItTXThXMVj8nbpt1IDhVBkPKAJNC
7G9qVwBX9WdzJJ8CejPwKBvEjmAfL+6XKM4X+adupGR1siRQYrLqr1/HS6YlMpsYl8VUoOAoNWp3
7Sz2myc79dHO3qq9ysfXcW5WquE7HjUi3yQetAsigQz7LgMFwYFpkvQkmO4mFYe1o6gt1yed/DP9
TvecwHoifrnMrJxp3Yy6Vxaf8VKMjY7T/4VPxNv7VCUfigrVWisFi+zR0eYJWZfPZy/tSKdoOKq2
+sZ+UxCJEIwP3cChKIh7g1RkTtP6vKvNENTRL3uWOroxro6P2i4NhqCUMFfV3V1n9VY7L0w/CiKy
f8WAhOI+UuMY3mvfAfrOgfV+NMnUMakiLwqfwq2Tc4a7fpSClK1Qo3hyk4LN/I3DLv/4FudNrgBl
sQTqoLOJ82AGmDf1rnf7CYkTG7rRQ2xV0HVGXPipgtjtF3G1ah4On0uTpXo1f3UwE6QsQUKO+AIT
N+z6eGpzln5daulQL87Dyjta2S2Bdpq9R0cadfbFftdNJI1FyfQu9CKspIuKjLb/9ERO1CbTRz95
ECSqixpFctNTAMR39o5mM75fElHM4KtG3J2v2sPE1X+BjBGfTb80GC2g/rrP35p2wxklEsKfxGmj
KhdXmtlmlg559K/ohuRrjcS/r5FbuFr8xTorT2hpzU5IoGDq57SDB0kC51Q44lgH6uLPCErixToG
Ty5C84EqB0sbhC++i421DSA/CQE6bGRpxK1pc4AM+mdSNSlTI3GBj1LuyXeTSTISWQ0MYqLO5N34
vC8IYugezMDmTzAwL1acxTtw1HZIWGetlR7gRCFfNrGllyOMiytLdFtrFn40IDhrThrzqawb/Ro4
m2wDZlqWMxGAvWLJpqiHcerVBMuDSiEOpByrEVoSAEUVYc/KJSCjiUK6H5losh29JyxcSKJek+2Y
c6kVsAsoEVOL7E6Hs8bjuJzCa8spGHciiMS2jdG3ckMGwdIyWz4BmlRnygKIXLRxdL9AWrMxy+4N
/cO1gLKi+f857OMQZovK1FCcOsFGaNfjduJ3raXp1WTs+5XvfzxalsMRhKGDIqmh+NTLtPlrXK8Y
oXYAhGHF09ookOfnMBB8NaM83SPjUrSiGzO87ieHBA3v1nKOWQ2R1Y2vAwS60jMlxAEr1Pza0HtD
UVE3omh0FXxB1JldOWFo9zT4R+Yu2E+VfTsIH/Fdk1JrdOi3AuducTLtRd02IFrLad8FoTi59g0V
kbkq9IGa4RaMkPygbd8xtCgOJrCGOM76yOw1quGQru/X+mOH0iFs4Q/Hv5HDvweir7zh/gZ9FPHL
l4eCU2LpCGnvUDF1TZX1JVenUfVvg5IPe35J9wBfVBso5s50B9jxIiigLJR8lAwwAJgavMZqaaCY
kVt5zAensaAwxMBvo/m3A+Wt+jSR06UqmiFGQPgRe6wPlGuilQfVK2TN3T/idPwo3GF477/7re6z
JTFBnIYEN+IHLtmRXTrKdq1V/PqTxuhPtHA9y+FhpaU5xusWUoOFZbOX0JF/hk2Pmg9Z8mzAvHem
AwdjqBUkxYPZrfLrKNx3A7RNYkFM0haw1WGx6IS23vuZfTwTl0vRY2xx/jwAOm1q2Vfax86QcWz6
DpwNyVFw4RvDFqPJoRzlpYD/e+4rdspyg9MqZIQygCeRAE8aHrayB5Pe6gz5uEvoSNY6ZQh7JNyg
DxOp9hG6BLYjmF8PunAyV7VqUAf7fKshqzTtQbfvaBsLrVxUW4WYsKbhskf0QCLA+1TDtJ4kdnQ8
thMO2ipGADyAb6xwqS5FGcn0rsmTOj+2uKt/Xaw2BLHuvlSngbywRLicr/ZkVJlzqLJmkdaV7Vtl
h1xQhxl+mD6D91QF7vAf6i3Lfw7kh5rgjsaEQSTGqPiqB2z+uuliqvRrxx+SgtiOjPYwyB/HzCo8
p485XjiIZQeZB1+ljt+ZJ5AhCBTuA0WjfzG93mtjYzBc3EiX4zolroOOCQq4aEnst7IKu9XWdRco
JxekMT1l+ulqTqPfmCFc/wJVGnyD1eT2PUUyzd9zXgnRcQftYtj2phrWiuo+9QjnXDHfMcMYiwRk
l/TWByzSZY+rxHQEmoSL1mRLQi5KsqBs21DUO2r4/zdRBM/Bezu5nH6FzVUnte/YAC5L59fxoNb7
dy17/EGitcWM2Xosf7J1cc9FnLfJAEZItsHtUyVrBxglKvANLMs1jkrZTTL9L0VbdW9zE6ofzP3R
0ZZZqHciUMWycY7+/pUNC5kz/12RZ5SQOcAvmJ2VBzzymrM6xac967MOFKm4incix2M454JcDSQj
hm2FHpwiom3OJST/1SArBooKKAxlptqKQnJewX9d1lGesQCTMNn7IDEpg9Nm5T+23GeMm3FLAmAt
QIRJgsDbzwM01Hxrm4nXEf0QPirMJT0PrCgzJ7MVY7LV8Ax1Z4Fb4en4UIB9MPosh4+MFvJuN+x/
zSuYyApztuiOYHJjAh6i/dN84tRFFtfdDpKYns2azoaxGJlrjDyI1DmhOlBOuN30onNQlFARoPDw
vZcy4kXW3dZE1igmE4G7ae6Nv+FEncLqjd8Jpdhp12hnlj0xOZ1Lm5j3FCQsBmq6zc5O50WIPrO+
9dQGS5PtgevjtZrGBLqKnmPV0aw6ZYHIxupE7cNp/fLaZ1ulBlZ6jtG6Qbaj6EQs7MvYWkFJ49/+
BOOeyUOh+g7S+JPTpcOiqysiEUJt+OOWagW8pMXakswD2bFAFch7FZrbZqg3638ocal91vXGqKM9
MfRGrbZ8vVOISbnIqMGosYEYqEielDvfJZGMm6Y2sdwtM4LuGNDrE6TjMzD7SICN+BijVCruPtS6
fS5q4ERHvUHoZCzUrsFA3hNCFkHMSSG0NGdwc8cUAwHn3TNZCZD2fbzOPGm4NYSwYJt7TpPTMUu4
r31Vor4Ky5+D58BFKg06EQMTzECCsktaXMkKLB0Hq04i+ACYaRxdIJDhxyyiz/zVDA5bmXZNg57o
lZvUOrhKpXaewAWpgiWfabzTU8BBb0IUf8Tvkq/wIsilRQYcpUpbvGKmyZJJWCROR32pZlzDFL2i
VTd/Ykzdzjei9ouQg5joWCR6E90aRSa0/yePIK6RVsyKufRPl44W9D6A6JJNOAsnGQLKYN/e2ahs
/P+TKeipl3yIsRvr+MIdLZKodDQEWFQVfReHnJYQuJ1ID/44tW0pqnxWb/RmlYdbKtbdgA71JkcK
GW4CmWMqJ7q9sRHVClqU8CXK4dZ/6LmnYlu+Y3OGA/Tc0HIBwVzXGfl38aT47mXMlIOKfp4jjttt
GNRDgUntbEsPhK/4YhkSFvoSPq8j5JmPRpfG0GbwKntw64rOFAQCYUIagAinuZ+tRDKWa99qQ3hf
lJ3+kddledEeK5uuA9OhQlB+vzibsEcu3XJccro4+6GzvQ18Iw3nwTxoNEAV82/LW9DYwBReMQF/
YjAWDlF/YQN0FFWz5aIa/zgEw28NV8o/ZEo6YLLiB4qrASYdTYT6UvDWesuwVPjAsS2yVG80fUF4
qJtzveLftZLws8FkA5rdlky8TBe+dnVkiCkCqDdPi58EIrKa8Nl7tWOPPKOD07UT1LbVo+HAOpzE
hrjWGI0bDA1AJEJe2COsy8V2/V6F7sVX3c4W0X9bol1Q9jfXMc1D+9LKxyOz2q+PezsTXX5PpgQe
1SlnlNaJU1L24UQV2aCV/4Va/DrSJCfiFE58zADierOxlh0wQ+w0iqf8u48DZS6vTpy0oYOzSMEx
+tjqXIxKIJXiFkRWG9n0fIBGSiGuVDx6Obp28EQTni8xGWSui8/2/9t+a3Bi/dZOOuikmBmq6zpe
pYI4MuIlksGyWNj+84D6GiTbr/7btlTbLyZwCshXIb2ob8kpnWRA1frys+GKYsQOhhVKZ1qa46d/
mAyYOwsDVf3Gjigxo+C1xL6l+76uPok/Hu8NaV2kPANdV3HcUYznrLCw0fJ2ep4khbWviaxr6B2d
kIiqU/8zxZOPxQOOk7RNxCisy5Snzk9vFHgSW13HVI7PFFX12+kg909Ym60rZmS6w+Tow99U159+
Vg00KAOnHJgszZ/GU6PPhV+nUxgNDSu6DLJ9cgelpF5hZ+r1SPIKdmzlaq3Tqs+JKq2plna3RfRK
LhWe2whOPoicAUz3RhBSHU+uemm1hT9YlSVl9iqu42eewt+OnlJ1rsuEnxbGBZgL18xo73VzHJ+m
W+7xQssoYoWcR/uZXoSjheKbOaYSZOlT/APRUM/l+Z4WTYv7iueK/5y0ue3zDSOdGL0QQQ0hxfXm
4pWaMeytc12FvZ1Byg/1MNXdRUUXsyTG0xuzVUGquGkAE5zA3OG44DF2nEEJDVLZt3RzBbxy1CLh
rLv8KCj4U6qEpoWf7qhKFcRV+HaLaKOByClbmA4/Z7O35lRD6CSpZ+Uv1dNVFFKpyK6kzeXv56vG
52UFXWG2EpLDMRro3dIB+2wkAn6uW/AEuqkMf6EERT+Ju4RD3ye11sqcaz/teCnMufKVXF5DxvU6
uYoalctb0arSqgpaPQUEG4v5+taN/c0fC6pcMuiu29tBW5U+pkMKTsh6UnRvtmiOgyNHMFQLtM+2
NyNKsXhQ7kHgfeX+B9/aeiITZwz9XDKtyBXGkiye6Kl6mdz4QVw2CosePoS0ieeAroewfttjaDZ+
8/g5Eb9jyQneGNpxU2qTau0dHT0qSNTQs3WMz9ovkzGPCLYJTHYlGVpbHILASUcywfba+KU04MuQ
6Kgs/Q+Dx7r+eMrTlfcNBoMOsO5uIwYoDv0YiBnGYES88PU3SGlp0VIJANdyDxE42mWGgzoB488t
EuHGvsw1CLDOQLRVHQbEbOZw9SQzoIMane8Y6thiE2vEdHEpfQj350WxWokhVxNPcWMGupgAZgLe
sotg2jlN9b1voYDC6OuT1woxJXicnAeL/fmyk91MoAOMy8HNWpqeYN1f8cNN6+vmVJGAtPzR1ba9
4M7OnG6i0VPo7r49RHs/6Y49LEU8Gv0eeIOpnWLJzCSBbTNrNcKXZcZdYWrWHNM6bXqFml1GvPzD
dYOtoytqLawO4hWo6iqHw3Vl/GTztZ3F2QA+C6G4S9HltPdDIZyvnwSOov2ZUYPO5AmeZHdqY5j/
I1vBGou19eAwbQqsMq8xLn6KRwvTuiZgzDR5MybLbpJOw72JLSuo1Osfa9LDc+QRyFAU1vTk8DZV
m/TWYNH+69izKvZbxhNj595R5O1KapMfdQG+Ww9fwGa5y4bLiACVzGL1sTfcEx922Oz2+RzW3w0a
5j5Ca2+ZYv4xkLyk/wGunjGdpM/ROZ05iz39Cdyu72sV+IuCIK6ebDgKokqkgFoqKZN5JL1YvNpb
CLnt1kWOUYx5MJi0+NkuN+F8ikkjTr/cI2el1rE/08/Sv9PXUfktPYnNIxSHjnIihzN+rVuDHe9+
wFEXtPcgImxETQB4KjlYSBa3BhyJNgX2L5Qpobn23iiYFLjiYxl6oSggLQ8/WVa4zSA6oF4P8iOg
YVReiO5ElKL85s0LEySSaA+/ot9IiAyQS4j8ATpHI40RDh+p1WmOEBm20tlGwsldJhfwkPpL9f9+
wgfppBQPhpFjlgcvvtjVmBk41EUiLqxyu/wiX54ly9Zgr5EVbHndp0huE+YdszDu+B0siLygd10w
5QD5pJ3SuGHPALkE7XQRW4KysUUBs2dJ3d/xu3F6txnGVp1sYvkfLrT4Tgq/JPgOmzIbszIHYwwA
SAa7Hy3G0cwPuKZ0Luoj/7788HzZ+Ety7pnd7ktd2T3sNemCKHrULBec1hmdCa7Twxleh3hPLyxc
+zDlaCs+eJbNiQn6Dyet/zVT+X4LgbHBsH1HNyK/lu9g+fprZFyuHUPwdUMG7NNGbK8Xqhut8i2x
/4vAoyMcDix53TaslUubE3ws0Ly5kOs5oM9/rYZfz2gEa/3vI90f4dDCRnxZEQaLx1O8jbS49LEK
W2azSb32MSy883kzGI/bchtUMWn/BoXMrlCZ4ZcIAK3oWhEhNbiTUcvPVfMEzUV4qct3jBm1IZBt
EMumf3b9GWtC44Sz7M51sa3kTH1CcUuJy5LWOwlLtMMGI3que1LWTAAQSutBWDDNSFRHIUrbwPuR
mS8YOEbs2GOjJZ3uozEdxzT/wWZ27lRcOfi+0obDT6LZKveWzS23USZM2krv1E41/mUAMYVrCTRg
RFosifmH5Ar55rYRfZsLT32zIXuU8vQpuuR/EMu+HpAztsNQiwROjx1JgEfRPH+btv2wsgheuY9g
g/rl9SWFOZY7l8E6MnA5XNvLf+t+cdPTofwEptQY9mEKqYltrRwMBPRNwSzLY05yD9RvZH6XIz/f
jPBZIhqvx+oWRsEzeB3Udio2mlMADUnSaR1SjkxR5y2y3ylecG0RFPwvGzuDsiHLehLl7OWY9VHy
ABqWhsQl5RdKos9U/OntbtUgockwR6KaixENr6jOXssYtO+HUXZf82Go2LEdvNJ9FDZ9dYPRFvAc
ZXDocAcKMHSpJmdsi05UMf1lK/OHCGsabH8wZD/oCl3R/crQAzjwCPycdFhAGrggjEJ5bZs5hSpA
7ya3gaoctYzksRXgYxv/dyIFCC5/PwGl4Ge3Da6o6t3qEGZkLCJnOBQ6b4xunEU+Ru02bOFE6zH/
iuF5uj+ENvg9uMqSPdJx51CiO063GuA3UV4F8shWtBZocmXtnqEJwA2lnUoRH4G+OgvPBUrbAyRf
OmwkhXnXtXcJXr4j143L3Wrp5eiqCc5xsID3GV7jRz3B2oxefro8pOtE8h/Z4Z6BwqEOv+bbQV//
TiBt36uTHW5lOtrxjpJvO+yzDG970IhbjKRdROf+5c+IGkmmNEFqRnV0/CqCD74GylEc3qCVVs9j
bGE0sIRYXJnZvK60WjS/am70zfsFvxS3W4lA52qgPVANgKVoquhY07GQooHCzHwtmlzKmqTYsKBT
LhnBuEE97KrFWvIIxJ7lcpbshRWhgJUnrIEdT6OcgEYDID7IxqiBkzc/20iK3nGlMw2zTQpi4pSW
FSZDmjiTUu/tSRSMX/UX/UE2pBsyRkDHEuoCnYr2ONFYpjog1/se1PtkJ+yIGSJozn10594rYM+T
+C874HweRtr/RMyKrmL4ceXXQgzbacVCCgOjLjL+VUm2+JKsQoJMy+1Vqmy9vDrCn74w0IRNLZae
1Cc1s8Qa9+uXpcT9dXl4K2pJUyQf/l8K19ET5fEG2GEXyLgTWvk5AOANAI6FFHGnKNp7JPkbECwj
3/+st7gcIn0Lfog0jVAZ4+bA0sudCsBLz0Txyl5zahDXTKJceifSxPyHqiWwc+XVnijPw+yrcX9k
bGxn+VX0Tnm9GAMUbewSmwNQpy3cFEgLKIw5CbM3ZkimbivKUVHznaw39cHrwSrC81hN2tV4h+rV
ZMjlCd7f0ZDZrx3XNDcHUR8drhPDpINPl0mrfnWkmZasQ1WQkfquhR1sSzdFV5qdEjDIy+9Pd/9Q
ek/wtRFTw+6HGu2/aDkEwt+0mlJqEMaTGKGvLiAv5Ua5GmsgODDlYslDXjp21V78P46giOsEYlNE
nNN/andBvLj94KFmY1PG6iBscQgovSIcofJ4UKIXvwjKKMzo32OW8J/unkGhuG0Qy5k2w1vUt3yd
RB5rulm2dJeWCOBXhp+fIgHHzq3O4rCJxsYd1vu2l/hj1DZsogZqiFtaBeZLceOrMb8QxqVW/bdz
UNlEBy7d3Pxi8eSwA43KMPAE+HvnaZ3xpXT6nkECsHtdFHQ5r/T3DKjBExYQxjE7R/9uUtSTq66Q
sdEA69OrV0np1IpW1+ul8b7r0FC6dMM8xfA3vrDOAIDuFIFwmOVNl5IVNVaJ5tz1Fk2w5lu2likI
wpky8VEj2rxFquLiUxTmokqzhVExof+Mf+KEQ3pwErTijHaWZazYj3en3NuGi7148tmcbPlkRpCI
LKCSodEWaUJ7qv9mVP/D/YAHqa5Bp2SA2OvEE6uqlZdTACmEljIxn8jIayQMkb8zy02hGM6eCv3J
ENo3XbRhoLPikxEGJuGWjJhV6Y0FlUFqSjQgVhJ3TXGgoaNH15bvQYGtIxWZj7ENm9gYaMCaosXI
BN2ITnWp87HAi+MG+hkPgeDpX0sWVIqfIxXjrYgKsv7lCGO05jiuMjo2xNvhr1cMT7VHo8LYxhH9
gThVHDC6mXXo6PosFFn5GZ80zUj8/cRtz4btr+4m+TT8BkwnO0w6q1/nadMwH188eFrS/N5gIeav
eEuqarbfF96dB6pqJOvdI+soHvhFG2gZQuOahPpBOxIsVNtZ5UDjC0xnWpJXbt/ABFu2ntBqo/UQ
FSs92eQWRS30PF3iwZfF/m3SwvxwE4ZabUYDCOg6PwrnnWmPdp79q8yox0+jhcU8e+/Aegmyjl1g
O/l+4JJ+SRwxEww3ZBXxJDuve0IAByjjGM6ghSuPuwDbMaaKDKXb9fx7Mq34SLCD6w7OX4YysgpS
D/kuQpqAVibo8zC+3B+bsnY2Ry7VANLeQ1xJakOo1NgYRSRnAmk1asQPIdNf6JSrqeThHSqiTq4S
+Go3Vy/6Yc8DSx8TuryqJs/CJlPWkxlzguT5KLZF6ec3mFcewz14HoOIf5hv76U9F7zxy2KgCTwP
6YZyIgCvz0Qo9XoAH0hlsKW1RVBqXRUb6y4Vj2uXv3IxJdYuNB+yX9vM5cF/eKI+Pwpi3yQ9VEUh
AK025tKq2RVA0LuDd75zeNfJrArqoGR8os6q2Ix3PZoxNM9wJPkkHmDkWsD6vcCXmgRimfD9Euuj
4hEvqaL4Ucmw1vbYbaT7qYnziEzGmeJxp6trAyJU6lGAGpUy6Bk1RIRk2ojk9SaRK/2PL58VRnJD
5z9r6irVfah1rYxOIWc5NGpOlmInOqgOg0iUowj6ZlF04XfQ3nSKWQw9GnQ2iNeSkz7ChI8ooPLq
oQvZ3fcoumOI1AIU58NCPzuLuUXWxqoADZAyWbg/RTqUuFTQB5Su1LKXClP4wu+lhmc1HWUBq0R8
r1uGE159K5qktsgtCqrP786iu5q/xR37srxb9w3qxVVzudpLvpwHFVwEIeg1HVewNx3b4lXcXLra
pcBnrHJtkv52QQCgMREzW0+VnKxbH9zElo7yyXXwcPPfQUcnHCO69UHFB6j3Mdca9Ysg4qCfoh6Q
S5t5Wuje7RFjHEf9+2/VMaXzACSfweZFzY7PbHNaBZg/q3MRnyJYv1Er0H/kTMgBNFdKyq2Yr25Y
U5q2ZLYNnf9A5pWvnDwuX7aGm3y+wBgFM0B5blzNSirx3SVJ9pBIqFEw5oYppkasGF7KQS/JGXxz
0Qydd5si/rR1I6sdgeqiqc1gyPBkmrbIizSVz7jF6s935diGs4bhexlZNWdsWgOqgDuZxtYKI1mw
mnooRpGSmVR+yLFcB8ZJWMtuL8/lWaUodArsdRYO2P4BeDMIhpb283m1TsZAqh/SEIApYxVtZyoP
mbbffGBlDHgNRRQ8XE61CRhXr8kQqzWFRWXAa1THOe3NyqoBE5gc36xKaVJt2Q4i4EdtShdOE6/R
xl6VIvy/GrlnYicSGNenKzdNjmzKjIUSkTCanMpjO7IdVrozBZ7EIFSorFriGgMKs6liuX0dctam
zMni6WTR16D/O/xjo9USM1wCwj+F4SgJopzAddb9tXgB/8aQxoKkUaf43b62uS0IqU/7ctaff4e6
l1+Qt2wi9x7GjqcRYr+EuknKA/UO8mK0aL/uvXjHMi7pvRzPkhJUvhzmxhsQAyhaEnmg5lhRFEJX
iukE8i/sH1MAeqUDo3zO6FFwvpkroskc97EJCoqskcGUk2OXboWTSDxykeOpRWtAJ+WzjyJm9wfl
9SF9haBor5+sgFLo7Z27DuhjmybUO7hi36e+vC8XKUxpUd3VR/fxn3gjFTzXwIDo/ADFy15CckcP
FZA8d3RlB69S9L0iYrNlu2YfjERrYqXfWR30yYEgrVkjyoGgb0O2IyVzPhIR1CWGgy3CnO6jWvCZ
dM8AH46upM6UM5ktCpn8lteMDCsMq080rd4rV10TC6J2jxeinD0TgBjq5w3C8FXd1etBGuetHrZf
wdVd6ieec0fu+e4hNowu4MVe01DD9chVLpepBV1uoUtX0GEHZvZPUvP5VcKxiDvKvDlyHy7msGbe
xGz/A8nsUIHIiIPgzG4G9U0SsxpR7tUtmmmP8Et+ScxI3GnxVmypY8nb/Hvo3Iq7qHMBVwqL1y1r
tVNOEXCMx60iSITccstsr9KFs2EO5xXuU6Tg9wQerdTNljGJ8lRUmZGomuh/sFJ16O0scJfD0U8v
qvWyFaJnkhckdLcv897g4g+YU1qxbvqOTpdQz8A68PCHLTSHeBXUQsBRUc5P/NfLkLQWzg9XzkFa
cT1CbOoAahh2rL6ZG3F6TpUZg2mcs0pxyaSrKu5owt77aufE8D1GVYOTFNybhCVp47dgRYqcuRad
IZNk84mIMBNzWRUKo+4diVkEnRsvthw07q91SkPOyIa+us0qYEKz3qIhm/Vp9I/UEWwneXwGfuGH
ro5miv4vBy+1VRfKUxD9llNT9+cJg/4/FyetpGyxiBJSPjLkEGXWF3WASUz7npNhCfmxVx4s+Cfl
1J50uL+NxyMVa/yWuB+TinkjAzwsPdy4lGAL4yFIyjRGhMRWZHaxuW5dBWjTXWFLmTPV4cjMkRxS
Gy4/K316G8vLT463S4KK3P2A9BHTYdgGnOUg3Sy1rmKrEMUESKP6dqpGHP4gLuQ01Kz6KQJh1heU
eaEsl9YuALyy5xyj1RNaM4ETEYpYRa0PK7qCOSlvMEmaaBY8r3Im98RIeYAQXb2NpQEZ4UMq9ttV
HvpjfJUekgsOuKa6Ld10J6wpaXD/Zdel/uN2C3/fqYBq7OaURVT8Ko5X2F36o/UtSsc7CJ0XTptS
vcLPpenW/+AHC4j0VX1r2eOmT60b+AZmVTKMQDWnJkqwqRUBgoTLX9O01QGJtJs8DQyd66OIWsZI
/r68qSwotXHSyiuAnidq2L+ZExbw3SiM+OfwNGRSOcc47nJHcJgrG19z1UHO35gVu+r5SFRJouP1
6zXXM7wADk8mINUIclJmdJX1Ut6YLfiOjzSwGNlBG7CdsHFY8KnPu3E1VEKNbBbC7i38KRuKwA10
WXlBO6eU0+2FrNHQeN6HIiyyQRIWF2RTKYEpvq00P/hL8HAyPGOP0iauWMoGHRwUs1r0NZVbrAD/
ThpQhLpARJaYjYYU2tiPlZLZ9CbrYFh0lH0F7lVBcCE74eUi5lyHlEO0m/Z4Jkn0nWKlmsINfUv4
G5g6ZFLXdGAnvEICANSzO0F1g8d42sBVIAgIaysKIt4aJDwLntUZ/KZZFVkUNHaCU7I0dqgBpmdA
OsX+wsMs8MkBCD8rZJZjAKfbBOH0KygKMtnrsN9XVDcl2fx1zerwdtBLmDcNrLq1P4T1JAlNWyZB
Jreu9CCiZ42Q4leaHXAzy5M8AthL/eVhOi/w9tUv/Eziv7dYXXmFMFbTppatdqKr6y9V8V7axilp
6gT7Q1wlc5wyTlhcZJ5iM/RCCz0MdQa3fVP9WD6ViS5J3ETKLdw+GMHb7iVNVBJIsV9OBMHP6ClI
4Jo9qiqfvfh2Kr8biwWSKDl8nr98py5mb/TvUxsv2/yjymWcTjpbjcPX19HGtgk3yfZOt9iiTko6
6+ZS8XHMGBiZaWr6r6lEFlCu1pdMLuRqCdVjBiooxhJR6jOQm19KhvO6qnpLof/pX2xS+OvRxcEh
z2iD3S9YE+kERgabpw297MSkms/RYmOB/XKr+VMCwV1MFYSU6FzbRVpHcyfl4nd7++aUFzm3rCtE
reBEi+SQpZqEO2/acDFOwZlSmhRI+3Ttw9vKQs4HxFY5w58HOeAf8Xno7oE4+jDBx0YnX75n2f21
LObJSqZZcH5d/5/Co1C+BK0WVL6AjXux+MxHUeCTUUVnrNmP+dntdlwwUzd6mqIdIKhXxm+YdBwl
Bwa5YrheV5MnvSXD38aMc5Xfrc/0VZJaBkoktmdJdhhD43N8Nj7klthQ7fp6nNQKA6/AHLtc0/+T
JKn+hNOhKGFHzFcYW0vmh3BpNuYeZoE9BvpqVK1X3H3n/2bAuOKN8/O+wdqFKPG6x7Zec9TqVC/c
rX1ULDH41GlSI+5ysnO5M7RnRucrUTEM2ZvXtuCtIfFskt06ktNudrd96CJfE3giG1LUGqDm1G+x
ZYreBxAIFCRKigCR4pRUjVYUpPT2OP6nriqW7OUa0d8Hb7GyiKqp7dAtsNwm8x6KwMo+P0m2ybMz
rGlAltS/+pJk1QVds/MFzi3RQ+Ke+pT3ZOsaa92IFTeAxUKE49E6BcOCvi90AeRlo1D2taSAmObj
Mwdp0A6qDxalppTMESrsI4WnVSPLxMTa5O3hEy36tX0124Q5WvoGw7XVf688m86D5AxnpklJomq2
6ntK53skaPl8cJxdGKYbAWbKfxPOQ0kzn50AD1W/CPIrjfeDseA9L0Kd7Ozvdkwckw4xsX7359F/
b813YZ1aZPxw9++1tw2rF4H1B9SQMs1cBb4ASiWJwEO1lH4u8M0d0PKzQ0T9J4YQ9mgCf7Ht9RXf
MU1DLDMIxenRufHxVHNINZyPLQXlTEVBTcg9SqmTQpsivVsngQ1YA6fkLOLMEeyfbmlNLOGPUFwQ
MZEQXcDcXGNK6ioqkNkXaGpHZzhASN5OpqWQyu6WLCf6PcOpWSChm84ajj7NoYj1gJJ4MKQWYN5n
IOXZyqCrCcWiJc3qTRa/M/Ce603z+T+rDcOakr07QEaJqZ/418eYuoKm1k/pmEN1ccFOWHYMwT8g
ewwN3OFjnpVddplX+Ged7NWycCQEMJz5gcbxhxWXQDZAlnAOOetG04/3lUkOfV/u0q5KUAfXE9gI
ofkYRVAGtbYPIQBle96UVfxS3K1rqnGsOsE2f9wMSVRUh7f5Xib0WAKWv1eB4gcmTdGC9xr7KzuH
0CNxyow80uVkJW3p9kHvCcLtW5mk1rxP3jQQDtnC1X+Dj/yZXuIjhS5Hq4JGd6o2OOr2tI+sDYmN
6HgOqTglFHHH1bHtpI3R6OFxteqrzcAQmOOVf0QEWacU1jQXTaNYCT3FNL2o7hL9r8DAmwjtE0Y+
6FejzOvV1Xp/DZO9PMO13dwNU48/xRdvRk07bjOdIB5zxEHFHxqc8j2mdslcX4vuMHgALmYH266C
rDWFDWShau1Xscs1ssugoeA/gHgG62Lec0Zhz75RCL4bkqtNbbKnh1TxNlhn6dbNcYmiL8M0Npj9
5SrdEq5udlx2WNShUjyVszNdVrjmTXiB4IDC0pZzpIGOgA6bTXsCHB5hJoMjrbGAGYJ7JBUUUufD
t8c6iKgs4v5KtRmuQrSbOF0mgR52pWqOFAiVDzBZQqCsvmkaAR+PhpZXU5jhFcvJX2SGFFXGhpBH
Penpxyp73eo0ayOsoeVBqqzSZWF2KDQ8CitU8FwStq5hbC5OuITPm2tG7iZiV2rZBzXcyUhAw1YM
w38T3GQU/oKd4k9cTtEnDJrzzrPWdGxk6JgKQoMazLm1mzy1OVilHmLU3d9iQsgcQdpMRUUZ+6hf
cM6DXnSQole2Uta75PZ4+Buq+AFnbK3P/dMBu6qiZdIbRt53wDJvzTNPqJoWClFZIRkvE1lhvXE5
NP87KrdoXQykbptrNqj6oxVB1BXJqwDW0vgvfPGfLGmdbFqVdRgpm12kc4feB8FwCz+XCRUYmIrw
76UvySmiboDChY7ziPofaicrKtCDCEiO7WWVIV9TgRTdTzMCVZpQMoofrF44XjZOVAWqzhqomqlN
F/fhlLMbHLi8guY7zEUSu5bDyz/1BFecAriT9BZHGTXOjLR3B0H/+Yg8N5EMlvq8LuV1Z+NwSGSb
jV0FQwHgLzg1RNDg+NZG2G0HItPLWJawS8dzhEIKRLT1pBLdroPQqVVmHTEeXjsYTjanpIdnPPiY
l2rRJD9573TznRGnLv5MyUeL70g0xIFvfFo+oes4i/HElQKSRCPREZHill657bCfab55PQoBQ8Dq
/NufqtTrer7AnGw9ob6lI5DcqMXFwdV1CKZanSOt8B78/UAHJ5vM/RsLWX1aYdPM7AY2kiFx57iA
6FnuTqIuhtWEoeU0qUyTpzgw9Dt9MU9Y1pUqgZY8xWURocnfinR4UUh/EiO2IMsMq2MVk5iM3kpn
a85kc8JpRwMc9LKiHpPk8mpLQfOpj10siq7AlfqugugoHVLXDMvvDYgsAz/MlzIpbt2kCkxBNffe
IUwhP/P0JuSNCzRG0zJHp8mEqBvfR9AvubUkrxxwC2o+xS8k2rx6GZWHPIMLaY0G/UQ3krdKpuHH
zjnpYYgFG/aKjC6RwelD/IlBb23gDMXev3bLCgLhL794hzegpJ1ZjPLhrnvq6fe0sbM6pnI5rwl1
44ALrjKbMptc6iVLYebq1fty9VTWJls9rodW7YBNhzpYLuXUleiUdDRaoqCldeS7bgoBn99JLst4
Nzxw+G3Errx3OAstneZ2cs5LAj3jchMAfoygBKOO6tELwgkUUrNPTDApOcapkhszDdGCUwVLGNQ1
PQ9GezKCwUUWepAx43k15mQ2GvjQ20sQub8Q4oPu2y/H0w07lcdOdPhDqGwL4gk8UqdZmmjtvoa3
QfsFC+M0BzKIijEOfZ5/QkIhbxMsYwYvfWLCRKyY97t59iVGU05ZeO4QAQYcfL5zACaAuo7pZ3KH
dFwhzsd2uqr70yeaOXxnDqWJ8q0Z42rCehte3SKlmPhaG+5XoIyG3tbiLlnNzMFI/cqRmT8HE1jo
qPuoNlJqDHI0ngOsVceyHovQ929yrdbID6TSrhOEm0b1mezHlZGVy3Lk14K00AL6xC+uFl5Ws0EG
JQgoL+qodrf+skbFiBBAaXm/O2U/6k+OYvAIhIgw0wnJtqAPWUiy4n3DVkcxIT4t4/IHL29+c7g+
CRfheOTQhO8NEUoW9otlNhAb85M+l6r2VQ2RL5KBN3PTp14DhaLWeR5CSzuP1g6XyFz8EhWRII6X
O0yPPLcYbuxynKT8sVN9Ou6peiGNQybkrpMZkoPXptMGOj+NZ8kSjDM1W2lgumsKqosqlJa+RKHN
+7jr9eYmWGbv638saqAd2ttIj+kDqFIgUif5r6qt3DYjKGjxBWYdbvZIIc0VaSuMvYTeo1gdT2uE
gI1egcGEbL3A+UuEiXHydnJtTO7j84bh5aFRU4X5GPZZKxzlia3bMWkJWKY2G7NytWHDiG3WzFwi
G5PFDjAf0gC0SQmd1iInLV0ZR19a2FDH8al28WAR/KHiC3SLTFxy9r1nMBiJilOFm4A+j5Mpuvr7
+j6dDm7cAw2zgObRTvKp5qf2DYMJJ5x5hy1WQ/OcTj6z8QDdT3hTOZRXgP4AwOOCT0z0y650f1ar
f7Clho3I+35oW5vIpx0/nI+k0Rq0jRd1EqS9780ZHYHwYBgJzvbU0p8tKx0c5j62KJoKksrSjelw
kSEwrDUGKEjPNHFl/KBt/8sPqo1gXb79D6MHhvyPfRkU9w7f/+cF/z+0EMRXGXWf/tUj7QzhoK/y
vtT8SBYXYjZbE5Tdl4IaCp+21yQEQT0jzlpNVoJ15D+vrHvF/GXTDYZGM/zw5nJs9iEZP4j+oo9N
mINuTQkEiY5gRGKw+O7nyolldNbIH7e2Tqs2xYzzFb0r+LaaxNcswCNJbFjkbXqbZmJZG1UU0ELk
9ayD2aBpD1Fm0ldENnO9iOElVSbJcA2+ruJCWDHFpZtiOzXIhZbHOa1iifc/1qBkvfEh0Q97H1V4
tPq6WtZESo0nVFKhR5x5kAcjCxtjxBCtq10Y5qScEX5CVD4Rn8vjBkEavHGzId2ZXNy6iUnV5mbY
DV5IGCL6dAKxO7RZTenorfjKZw5AVfbg6jB+Nqrt8nWS9quCpmOS9BgvCkEyNh5s7wyjlsk9DWO7
uNxVJOtfOEYvqbh/J+xxb48AffBR7zBTPRx+KfId+boeWt1+Inkla6QGXcfjDS6Qf1BUiyZ0YQaR
rvWHiKmb5Zii8UrBkMfO+KGGE0sheJOKrRfR2q5xL+5zkIAZkuSTcKk8bYhkFSkAucNe84xMtt6l
ZCihUct6Scgg9avaG2CmeKDksbTGE1xyXpRiUKvV3T53qytY+Fp24n+0b9Fy2rLZTmMT3wRq8/9g
Kpx8UOKlBY77YrBlm+asCfk77ZbS0zeiX6LQy1lB7PrMFI6uhCIGVlmmnqbcAKI4zK98AiLa91kn
y+ptZaoHqdTQcXLNGh2R0Hlv3+9AyfuH5FKrPU8Y2TZJLVx0vM8fSmZRB0FXsmoe+Mbv55px1lID
6bg34IsHehG0FsxahRAiPPPz9JAmi/PIHeGj1IQzM55rwDiG7JQHsdvLPZXJ7EL1qn8TxuKRE4uD
tcIWZOwUfkSTCnUlyOwyHRWfsvXGxtrxs6Obhb+Y9IK0QVrXpZ22NenoDwgRJEA/fcSEV/dC9l84
qUdiRu/rpJeVLs/axqoBiuYb2atW79cMhaRtm2krhFkQYxVPTtFHMqPIzMCkJbwdS5S3ugF2TO+L
KH3WnmbEp0+1Ku0/lrMyoBH3tgNNTXeQi3FlNrVvWtLsY0dIfq8IJ08t9UDAQNi0eCkyXX39Orxo
mSSx1Ipp4JQbB2H78ij0glADMoczEqaZyLnm3DLX40JLCmc2AoktzGrVCFKTdN9rnbyGwMMB1T6/
acb8KRE0yBW8ZnL8b2gMmW/rG6PZ3hw9sQBEt27avDX56Y2b4qJPnDlbRLif6wiAtkTKyEQcSrBQ
zhmxhEgaLIZhE4ByAyLowDG+qAppXri3TKqe1uxMlqtS5WHuwqLquUAfv/YPTFgWz+ioMUzOS81r
rd1Jy95LvLlbQ89vEAAF5jpG04leS4cLoZ+nlrcnlRZmy3/ei+Ga4ZFp4yCDPZJaqgwK4C9rg1po
k2PONOE8bMo9Pde9rIN/+56h/fQfqrRiDWx1h6wi2c5kDbXXFKFXAjQfJOzU3tGKOGCFydHUna7s
ZdOIRg+OeFrjeYqXMgFsnOqH2cHTKG5KYwrlJHLxN2dU8l/YeZC3pHSccsVjAsDmguf7yQ0fjGYp
UuG+i2XTUokI6gO09OObpM563DdBr2r7g6xgTj6zWfaMnGOn0vL87lRPSq0alDJxaaks0G8JGKSo
75H7e4A8qcolx76X1cV4nbOfKK0dFHEEiAoL2B2hssqewqB4626u00XAXOiM0vaIXDvNRKeb1wOO
vooyWQUouZRFOUA0z8ilaiYeGYKkyHAnc87jTU5V0pBhqZnXcaU6depLUPyQ992G9NZ0NZWHSlGK
EsLqBGuVmC6YziY9KR5ko07WK8BJ7IwM++VEFnTqAkupLc5F1EZOKnqg6d0v5TTt/AnwAEUJrGmV
yOqgJoCkw/U2fVhgyJ64bqGiwa2zULqXQKgv0GpdsLJ1KqAi50NweHN1z3q+1tujp5xf1s6jvsPJ
4gtNfPrVbUCRnMlPR99BXhEKggT6fxQvyDKfHw6CwPRjv/BbjWaEQbmo6POC+eZrCRDs0aIeVjWH
fPP3uGi9DBvJRuexZYNEaBE3GHbALxUGVldLC6qZ44/CqpLNl9YJ2lu3e5C03Hg4j4BhMKtoifns
TFv1BDbmTRlPw4L1r9ye7mT1ZQxzU69ZqPoJ08kDEtsuBI+W5CTYF/4nBlD65H+4hNAYxkKaFJ2y
wfnhdnB0TuTOTucE8GxUFHmZm45ZyGJTB55rlzWIUAQWMBm0ntvmDItag3w6+M4NeEmMJxjRvQJf
QLSjHwokW/97hcpTOw8JuxuNztHCxO896ynT2Yz/Rfy6u8vZenDAWdM5Dw0GqJMHacEyH+k+jHD8
0hurAsHy2xmyYoAhQvCaaDzYfYXXKzFoO09uKPWNm8MnCUWpfRpEPORkogrJ07+nHbD/DHfD5p9V
+3RNesxi4a+VeKCqXx7Ca2xpij97Y0/O9Ue1hRQyijSuwAPx5KJ0CVDBGVWTiRV6MwaiCa+R+pU0
L/RxeZqzBV1mOm417MwLi+aGW6VvvPAjfhDRHRl0pdvAl4clVyZSExKHczJtl7XxFybypvnnooV1
q9MwadssN5G1EdNSBe4dNc/jBq4Ol++X6Bds7+TUGFCrw87fBCW6gF1CdcjbcdCIox1gnCpCy9aR
Pkj20Fp2wyuunqthqu2EMVM1v/ByRnZn8Ynmvqb7NTHl1CdYLuOto27+16tqVYD79pX+sAnwNCuT
vpSi6dypymEI4Bz+jGjZaO0jehJ6raTrDuR/LpB9RsnQlBfDbc4GoUmn7BmBjogC30LbAgTbi1b+
Ekux2Mks2isNNNsi7kmAP0GmaHeLOs3qdLWkwh4ODkh5vzrRUcnD5bGnXyk9gvKgQc6i8bP7BNsR
uC9LZ8CXt+YDH/J8WitwRJnj94Y4NeCcohE+96DbMk16dqh8BRq1XiPyv98IvfNxjI5nje1eUCOO
130jOsaVVkdl6tDiK2P3hkUJCJ6IWPMQ7xn1BcYvRf/uCZ3/q9BTTz27zOua+/rB8NBoOXUeCrvN
GO1P+CQUZdmHzFr8EutwOoCBH9td+3fpeRRpIXMpHNq0GJCSKRxokfFUcqrXiosi41aZVxngUDXv
rYdy4nYtzby+MzgBovVf0NkrfKkiSH5nMpMNdhh3rXfi/gQPRk+wa30z+jFOABZP/NSWVNyAJS7g
CrofQ9kxxjtpBr2TUm/39EnGe5SYlRuGBFH5/f2lZubrR9jmK6GKPK/j7MfkVN/xSxjsxburwXYU
+BD85tsnkD+db8v2vfh4+TDVVBtUrXIGxJdzA6wAO34WwnXc2C8Vych92+Hvh3/ZhNmn7jePGzXw
lv6Mcl3pYKkKE1NxutMgyOQTWVuDkYhQuGkTQu+mA6zxRwY3Scx4yFDYe5WRysd2KanlFITDHQwQ
c8qadhKV/b3atVut+zeSpwVx0r/APiCPvx3Tu/8qGoX9EY4MY+4kLW8gaNSFaR16D+SnsFAVtnwu
MxsvPT4UVck2EkgQU2Qggq9ljF2Z4Kqm4iSEZOo5SF8E7Xza1CMtoUElUd8J0cFSYoNQBQlOsDnt
LNdz5hyJi56O/9wVBjtT9tAS+bg2eRkV5ShrHzK2M186f6LW3ay91ne62L3oTm3GK9Ben9A2D144
sAqwTc9qZz33lPm6rIDNh1L6NL1W3P+K01ZXAlTh84PmWCabuajl29JYw5gLD6UIas1wOEhCXLBU
2Xz2aIbeoNb7ufg7kuUc9HmoIDqYTeCmEKtfCtylkVOUgvCACZmFJZdWRjr7LzHkR1XY7njJUU21
vLJ9oVYuhSzS9KXySaonPDPeiwZ12C67AITNcXZlbGa6kV+W37ll9DHAsJzJ3l7vYRyCtCY9dWMm
GE/Htxsfks1Fw0mryPrxLkVHMaYrMiI7SnrKzNKjuIGHASkmL6IGZIXb43kWvJm0CzR/bm1jfot9
RG75tnYalNnLLSVG1juBj/7ljsJYipCdKx+g+gmswk63NlfkVeH+ojKitzACafvB6/r7d7fCnBeD
cm4i+qGBQLuhnr7s9fd5RTmPxxUG9447j1Nzaq3YlbrKUxCyAIGMZHDd8tNxXq4tmNEZaTWW5fTI
IYumIUAGopN9DIzYQk4qzlYJnzGeqiZlR3EZDRR6ZaF3qmc9853L5js7YsVaYkPs0OVM/KP8TR+Y
h/8OOBwNl6eo3LV8B7i6aDJ4WSJUZNr49e015sZCwm66US/tFN05w9eEMm18Svww4t2H1pUYc0FD
QDGxjn2jCO5mRj9upxnBzzp884EHzVu5SBnMCWCKe2ls2dZvVm4N1EECnFatgifiOz8XZzYmSVMy
tQHqn77+15K8PCq6a66GcKSZasaSxmT23o8ItWwheFnCUb9zOVtB3WEH0ABJHCxfe0Wwba9Ep5n3
FRdupB0QDnBPnLUuwoUSlX3JACzplYQwCqwAGmuIo7zhBsmG8HE9CD/pXNrzHQwkSrohqC4R0gfR
O1hbDnU3XwmrZt1NjMx34J81Mi7lfdKg3pNiFrUYBDylgtiJIhhcK2VgQviGs/rXaft7TaaSjjlo
7cIhfQ+adZe+p4akBs6h/HPjs1Keo5bdYy5KoWwFwz7CCP5AonjpMQB0MM8zQuf3UASqMGTcugAl
L4jtA73BbwRBn5XRJwQiE+WGePuvRl9PgSCuizIQIF3V3d7lBPLaHduHYxmy5VMoZfoMzGFBdf//
NADXSba2r2QWOJS/RkeQsqP89bjWuudS8mSizymsjimNnblTkI7WnfxaOj3nWJW8mmWmGeJvyu2s
4o+FmkqrjUKIGNCnJI3tgoH+fogx9jFhFfs7h3mzxdpSb52QCZxRAW0RvMxal9AKm62MbH0cXZL1
wuP6YS30YzG6Hg79WZNwvAGKgNRFoA45beTfN6fJI4+A+E7031sST4Zy9CaPWm+NsjPcAPy4t/Ql
M2jSue6V6LBrR4uKTQsCWOorI7pIO9f2Sq51SfV8eFOfTyKuXtTEcRvNJDRSnEB/qzldiDUaTnad
d7/6yRDZnhD1TOPuPyNIJDcrlu/KBzKu+VjZjYg3GxIUpvYeKjQEa2eUT+CvNR3GctrWGDKR0Bmc
xXoWOIOlp4WBNYKxltoJ/53SC2vEpvGN4UlTP9d+lJTO2J3MUS2tU/rzHPzTwy45Dwy6ZFanNTcd
6wSjDj0MFsSiFqrQznzXORE8hLsX2h1QsVSju8iBo3iXBl3zmom4hPt4WWgtqsOHENxB2cz2m+tn
S0nUGVrTJtgS2S4V6ofV8v7+FJDCOT2SOs6PnjeOU80saSlX7hLVh1yJ0MN6j3nWPxthb3fPlEoR
NFSCZO58PfauVy3VIPWWIVmS3PegfUZLCjd9MNopdEj2M4ctyqxAGhSbkz20uhd8IeIJ1I9GUhEh
39ZM3ge/2mAVoopakWiIq1bWxJ44oKWVvo59mXylpnIzICxwfH6aUTLOicx2T1Tns5WRmWG1DdpM
LCC11sqwFerkXirzWxQcujuZ8WCAUAyfvTzN/KNSemtg86VhAQQ2oIqb55rjIMiwDf7BbLMAq1TK
2WJvFfWdayDdtYKTnZxpLMPzZv5niZTXWXodkzETf7eu/839V5mr7M8u3fdcaM2Dn7Plng4CS74w
p8UyCYT16uDfkFMNJi/XEV/NiKyV3Vg2oZRNshQU6cIOUQA4judunbdToZCZxXapxQNqIs4GVXjR
r9bFrZGAPLLst3dqEHcInKi7RzTE/++0V9gepeGCYcwyUX9kfMWMOSt+xVIiQtNbaYkQG0fYrvT5
p7mn65xYltfbK4JxTv+RwWJNu8VQNQxyFpDAW20ELxd7LvnI1RDqSROzYdsXY0q7suG3JS3D70Xn
gC9LAQsP76OSmPtmh0t9RaZJvetgQ4VMSNeWSZzsyN79hb/i4YJ5AwnSVvs/0RHwPlF37vL59ude
ibvoU9P5CIc/KAmbVcJiWvyftGxKsWCjReH9ddxEZ4maF4E2m28jhE9MEHjcaPvRqphCNNqfhyKh
MYvDupClkzo/aIe3usXW0ySdGxsYbZ5T1N6OjAnlKNvevgt34bBNQs4DpVOufEL77E9omIXwD/sv
RmA+YXhmbSfb7iFtzjnOy2+7Ry1QFRIUd88cCp2M7ubd56DvPAlLGxbNgHwJx7aBWubS3Mn92NSb
QidXxxOUdZ6Tg4lgAZsisuyGOowN2CV1U67415F3Oevk+oJ9djqN6MCRJANuYg2u9LA4lWRQxi9m
kdNTv0bc0k4MTneYuOyuXcL9lfxaRGbC/h4K396vFcGnujSI0dv1k3J75uWdJyEMZDbXRyBVqh0T
se+eu3Lk5RxxsGkOBDExfYn60xygt6EW1RhlW3ct2ywtgOpxJhDgI0f5TpFjfquGYQdvwdyf6tjK
BlAudEU+SbLJWiXKggMwhvQNNufittDT8CUs6J8JhC9WCTtrUNOu5SINrZL1J4TJ7TF1eH0mUcPn
n4cvBzf5fSI3SJB+YLe32HkfyXWsmSbDRMyLKZQSqB/KjPM7aGnjQX7vbHQCgtmWfpfcWqI+uZod
3kedUiRdxYCgWUKS9kFrCGwOzknTgmR2+Q0OlqytCD9NoLP3qzz7pDeX3QwXxOKy7npvlaEN2teW
0CStbRx9aGGnTCYunhj9k3HCzHfzdBQVSryshl3bYEb5MKeqvzTGYPo1X53PuO23YYWGy2pVsiSw
9+4+LvVGipdGiL2tRteT9e3ktBg1V3ziOSHb1drWqcB7I4dbZWx9JstDgjRf5gQiUZfEKC0+Qcm0
/UJKIEGug4J/ri31lYp/l0jF8q6txCkFyfMgkJMNlHHbyZvAg2Em+Tuf4rkKCxYiZWYjmAdu4pPz
KJ2+kxxAoEzp/ykFf/dhx2moDY6KggLJsFWWnZK+W226Bh7TJf6b3HPqMB+QgRJfzoFeaTd0wHsp
v2MBABsBf2BXEIXeam0/9zdd2xrZd6co0LLGoFbqCGDRVt5qBIlV4AfIXizv0ZcxBkNP7ZNV0cDh
pOaOO6x/VFgh0c0adrpYTOdVg70fNXQbs6u+wtzQ6a1bjioikE1Jo4RgG4GXRiIP4vkIxMOB3SWz
N8DFqNGCTusts/B4uz5EgAdm84fV3mXhA5Ew6yqunGxYPnQsuy5jBe1Gp8UPMYwnUuIqf8YnOV3V
9FBBgOEZ6S8L3M/lfG5OXDSpeRAo5e5ddWE6lKw+g+qX8fG9eiTEo5MeuzznRb7ZZb+CtVf9r76r
CNWHPCIcCHu8raRgpt+Uyj8ovGrf9Af6+ZRqVIVcxRGnaJZ/abj4+GbfQXbNnboqOkyxPZ9nJhve
80V9VNE3b9YUYNaS9ZaugxlQihsltyM+8iEWVJm3d6+9n5+UeikoV5fmqMYYwXCO1Q9afo/d60Fv
hb2rajcI4/GAy0bZjS9kSQuMiuCRwybLPWBOIAhIpaOCq5kSl3TgBva7zW+3eNSwMIuP6Sqqq5RL
EVl4igXDAIkOxobhdH2jynxVex3wchLUeHB2Xll9S4SMNMj3q7uUQxOUfOVRQ7bogCQQKwZaJvNM
rKWzUB3af1psa6/IE4ebXOSYcNT3CbXk8cFkAQ4SAzZIu5ycEPQ9Czzm/m7ZmlHvWI6JX1bcwm5g
40zIUJpmiFWnIN8ugWXWmAaJe35irxD/MdAEEJWbTIaK+EITY4r0p+eeqMGku4KSXkxdrRZjr8Ym
XXykVfVmccHmjNJT/hLw2Pv72I1RqMdqr8psWg1bO1bN5VFHxknKuT/Ab903SlNKbsPege0tcz4o
F+GOnaZXkUdMKD8/wlaq5hWZ3mXk4p9Zx89Jbymgf0fF0EGwOot+o7VRbG4KWtGNZnIz6jmFFLS7
5b6U2fXZzPX0+FQlHo+Pm2t3foyTjHEmkKsm3dc+1R8IGQRzPw6dDgUqbHGAap9gQTZwjDTca9lr
xP1mC5fBFFwF9Ucgc4r7ekZNqv9zNdylty50+j9kjfB/Bk0+oDiAtYVkVfledub42Os8ousqWZzf
+JO3S3qzuIx0jWfVLZu+V4HEPTETJcc/cUC3ZDh3XsqxEjq22c7KicY9UtV2/uGAHvSiPDg8Nsnj
vz5WC/yJ8XNrRsN0pkdKaHGrF3QijyMLrb1v9ArKfZpDDLbXj7vyfC+/163rCElW7qLniJmk9/li
YvlG3m+rO1X5JXWfs+xpjaRs9MOIIz1NlBY3dzmV8fO8Um/qYjeaz5YNh74ypURhhRoxsuFbOM+7
I1iOTgUK0RvjI8jAG3iWF10KtRJgRKj+OfDLRiQ5FtEX8u/CTdMMfkv096mgHQ3qBWMMcgCPSAWG
aLxe44UweVP9nR6f8r3UdCoQxYieUgVhZ15zFFaLqSbSKgnuBgV+B6LngYBSQVuq+A0LA0XTGoqO
p1P8nPO4u5u+PpVBkj7MsYGLszsRpugnJec5/PlnqsiQWkZocFHWWcSzr/hQf7gBMMPE2reDpujL
myelA9EUDcZgIuKm9LJtiOCGKhEG2qxXtLzXTbvQrtdCYZE9hCw6k78yolQpbj9Miw36hHsEsh+Z
88K0XsO/gzHqHkvRpc4Zh1Xfvg2W5mZitWl8WU0+Ncfe5rMkI9dS9bRmNIv6zhzOqd+3BZoIBUQF
n8BWFROcsVlFuboZtcvMNzvcp1WpT+OG0ped5K9KYr1YUDDMUCZLATdxblDQ+CSnV3Pu2kbz09RD
dKKlDARvylV4I2n0g5r+Egab8yGgRcpy5F+O0zQyhvRmyyMHA1mNxKnbR4bHgj6+p1444tVM0iJO
swpOCKhmYFuhzUeFbzCKmSlQ8Lb4yj61tBNl1j0uULEME1FsTu0EACxpMJVJi6X/DGOJFijEne1P
FqThmHoVFLsCkLOKf5qt//bhMOP/s1Cb28QV3nylUu8Nbp2+A+/72sJgBsPP91/EqzoDUGmYQq7+
HmBFrpAiRmYAK03S5cxdGY89DUk5xP0zCUFKNnha+B19L74tsal1HiIniUcRF4xVXxzjt6Kj+zb2
19Z+jdmYrjudxfLcX7IZ9Gq9ite5yiUO2kzeOUTDg045IPR0GVi//EZeKAUTd3/vZEXEmQlqiR64
bIsAzHh8L5zNjpXjCqLXtcDpWI3Evee9umt89iQMXGKIDD20sn+vc+tHCb4RcW1KlIQhbNgvR14X
tpOEmfn5E39vU0YKPzG2azoWbrhGUtdR0JLWPnTuTrbiHaEZM6lEaZz+6HkXQWDg4qnjZr2KPDkc
nGanAy3Q8oKYB1lW/yq8h/ATISPSP/I8dfy5CFfwxtmi2V5iptQZX7hzfOhT/+5R9WB0EkfvMz+B
d1IXhlvaaUm0Ztm2bVJOd/GN7+3jFh+polOV+bZazZpAdp5YfeFZSz5neTmbh3BXpEUJVH0gNe56
Sy/8f8uSv0+l1j7SmTws0iDbWTYXmaFiZLUCGTx72UHCN/ijTtIDqFpjI+seBuNb8ljaFecZIVm9
uo+gzAARR2bwoRosAIe8NinYFYTrm/GXRj5sudYO8ZYQh9Rl5Iv8XAuk7xwK+P+zGq8tuBflxbuo
PiGfSwTnNYy/D1TfUsbTkF8nChE9TlPxTqrXHahxd62ea189RcomzZ0VP2C4Hxwrum1fGU5w8Kco
VjtRPu6tG7lSlK71IX42wd+FEkxLFYfKBATh4rJar0zvEBDBbZmQoBv1+VablhE2c1XXaoUh/8Ns
G7Lvum/2OTrqADDb9J404djDRBtFMe/49P812LZcfHB8vVWZlooqR6L6SNLID9O9x0hNhmJ32BkD
YZ71Qssg/N6otQUlTzXzRhLJ6b+fFHIjBXe3pElmbsxGNyguQ+aLzla05ZHLG1jqhy7Q/QOqgPM6
NMzVEPqUPBE4dVTLcEuoYOfUX1ft88Uh+thhNTbZCGcAvncpZ9JkfmASGkdscl0EPFhWcA10l+cq
YSDzabU3iKvSOezVth+RG+TfS/li70hOZ516yY+nxcHBlBQc9Z1r/lfzG4nn8PiDhbvvBU+Ff7QD
P6iSGjMaGeRNdGhB+t051dOZEWzatqgh/1xGGNJVuZevMgox4mGcxbLs+lFxa9rZRYvuqlEpkFW9
K2B8ib93uFvDRMiPjtifUTGbCKvIqGdp85+hR5Z9Y7uN7yyYkASkCgkEkw7m5nusD+tt1d4w8NUW
5OqPLa9AI67uhYj66nYiOw23LHY8I+2mkZ6GHNEnwTWK+GK6KzbRy5WaLEJSmsynldLqDCUwAhpN
760PBNO0ub/5FihFGqi+55q6s/T1OR1GDl6LdoZEYeVtBsM66pl19MfWunA9ur6g8I5fFrgotFjL
S9F2sJaeQKxW4ehM1b+18AgTojnyEOXZVqTS05vIxqoFw/9rTh7pZcvNAQx0/UwaJFCg52l8j034
fK9QNj1BftBvdu3VXYG9ziQslTPpDmEHuJoYR9O+2ijiC2DsdoO1SipdgbIeBChbxRl5nU4PyFed
rn/bFrRNSDGT05AN2Up4hp2jLim7Risa8wCPt4n7mJd56BlpzTQof774kS+Yujzv5Ji60eiNl0IW
WNp6Ucf55ov0eRP3UxmW2FGXTMLYB//uP6P71+ol0bqVQvsnlFMHye2w1SAyFL0RovOqQh93KN90
Lcv/Y55DYSLc+cxjScv/GFvXgn6fhLtqPCgPveO7o8Uo20K4ZyzfdSLbL+3Z3Pmwd4yQOqdLuhAH
P6chZ7QkmScU8ybNXLihSiczJ29QjK80BmWSN48XY33LwvfbD9BfEHwdRG+vUhgJntA6lGl2iNBB
1LHp3zIAaVc9MMGLkpomT95xBPR4v72f1jU3ThCkxv8ojgFDNTdN4LNGAsuRiM0GvJ1FdySFE83L
FD8KE2giZ0HveyjSMG4Ow3/plxyrxK6Uolf0q6Vg2QoWqVmU/1kydTiyDdcuA7ZlBNaNyFxE9B62
Hskf9UVRhIxegUWfxDLVCzI2w8GJtdJ/5U15XgBUvyHr+q+mSUJftbgL+zp+KC/z2ama1EkDN+Hg
De2msily6WvgG0RXAcNmhzsTCrmtVro0PwRKzfAIHRgoSuw4cNnLqqrGZXy5FiosiYgKx857JlPv
c5l7629TKinUEcsnAXjX7eZwPCvf4kkquTwzKL4O7DZb7yyngKOJTGZTXLuaTWcjYO/Ss57+/tqS
wWYZ8860ouukZkvE0y0YFb5hzgpDzaOaIUibIqP511K7k6aeBHGksexdwfRBGXGSu8VTSty46npc
JTOo25upGEhxI3jtxRSk3tG2ISGnqoxTEHddLJE2Ds7oe3X/zcUOU9ucunS2IDa2/Rt7YbTR10xV
4oK86jd7IN4St+fgEHjztjxYq00YuP2SSsWz652nmPE35phqBDwo+n8YumXcSkv4ef5AJe9SfIvT
msUonQPmTkR9JkqD7UEKlN+wtRrCmBNSlHIwgFA6M3IoXOdK+suTENV1nQgWJw+KYlqCgNKb8/XI
GoBxZcrmOiLkHGGyltE9yA1PqEZjgZ9O17apR3LKtRsZySS2SMGvFJ1C+J0mkA6KNVXcZEnSdzz2
nKYjH9ZUWUDdd89kYAsssUy26ngSewHoANlhwGxFlCGejHdM58UXFK0+CMn4Kl0luMWeJf+UU6I7
wI6NSZCaIP4GO0PHpdnLY4c4GtCtskLdWwMBDQwqBZX5bpEEeY37NcFT60QFoEO5CNSpW/Gntczr
hoZifezNrvYa27PW+oILtyrhfN+SC9zWJ+Jqj0vYYjD+70/kW7jvPHNRY8KIw6jT3EuKUG4r4Nax
JBo44f0RubdbZFziEFz8vnD8hRglRFdP1HcvQdh0bsV/6GpdwBQg7fH0g8jRgH4KQQqwrSU4pmKF
cejnjoG+79Hwd1KkSfuYma6+hwlEh2Zd2lwNo9y/upBlcrQX+tO7C/YiBaVc7tvFCkZRSnBVhsmp
nQ7Uxz22qmb6hQosIILE5PA5w+efQ3C2Hhx3f42NISNTQhdbKAO9dMCDwBMjceeyK6QQTWwhhY+i
TxQaaA201qrIwboxRJgi8cKyRZCIeMPeQsgSpNjoC59Qq6ImtURUxDZUiuV09s3424ABvntdRGxu
c3H2R677Z1sk8wDlV6Tb5rV7nPJjtSRI9gr7agRUprN/Ohw8r9/+tBRaeogkjCldANxxi7R/gZce
m3RLmsefSP/41QnaQMYU0OPlbarzida6a4ZhkQcKpMXDp2UrIW7HWHOUxUtcWhMAk5U/MHZBsqtB
fe8XOkgVW7tWdg6hjhp/5CnLOKjy8GDP7zi+IkTXGKU8J1udLB3/kaNwaZp+v5AnBtD2NHxiIxo4
mrR+fG/K9wK3+zLjC6Y87AC35aBkTdir2kXyq5Fkdi9pC+epZQaGBkQU/2EQbw/ZskFsjZ+MWquy
eNTji+NHFoKyiyvGDaDZ4h5K/vZlfrLH9TMu/ZCwsJpt0CNUerhc/l3o7kDU7P9KcsGPdvP+sK/O
cif1mKEMb9cTNZx+QlnTi2agzYUdfSEbVzrs6eR1DvGiRbg7aK/4Ai1LM0vba2fFi2pZPVRYnZcX
+UFxdx2aYKDJ0Qa+WrWqs2SOEOvaVJ8ETpB8XhtUDeuEUJl511OQ0DdP/N6dOQVVdYdNWMEY2rRG
7nhxXCrx0pNuRoElwcBxaFGRze/WC/eZwwFv/7EoIa03WU3B43OgB60+06R1MW79OVgO4GGMqupc
gZwH2PrqAHtPdgyQJfydHOB2Y8o+NWRxYrFw9zJpJRBTOGTbWcmEv0EGvbw4wxTvGpLpmqb9/02g
i+UkF7W/KlYgaLiCErxuSIA2z3AS5vOFWIpclFtR5ja8yXy9R3TRBqn5H0bBbyfOJkvprh0bbkfo
wASVZevN3Km7zWxXRBAFnl+t7YcAIRAVo4yvPCh1q7mivyn1ypN47ljju9NlcBR8alrFoOty8FV8
iP21vROFFFEWeIjONRvsEzkaaSRQmQdP8zMqs5m64UARRZkNKS1nBr8vgGSooVzTBpHHo6dSuFiN
/p9VvyImZZew9IVQidugqU0XnBZbGJD9Rr1L8HBwLfRgWWdL8GDZ7zm0GIQz3S0Wv7Pm2/Ty8ndb
tMySE6K17ite7HYuiq2fRI9jP6noFzpEBpUIvpwlLksg5L9VzERmMN0xG7xrL8D/vH4/UOyDnoSp
t6eEUwjR9kC3FXMEM1HB59G/R1jy6UDm9kLHXl2bLOQoiR4sujaYCBlg1MquItUIVk+bVfrOjUNW
M+5VtieUEYmlDwmzy/prM5lw/KvVBzi1rCU8eGAKLCM4kRtWHVdYCh6lKHQ5kXurR3bOHOmjUt7c
Rek71CCQxQjrX6zz8BEm9p1H47/54pIHOMyJzczo/wOgS7sIbWV1mioEocRkfLoXOLyI3RzSQqOC
K3nh+kros0H7PSivkJLX0PNl2HvuyHh/uRyukb88oVO4aAU/j44n2bSAoNOTZqsBMh96RjPdBCtI
TrwE4oFHdZwKeh1RK/i01FeOzk4eTuCKbGzw6LS34FDYLWODhmaQ+Qb3omUl8nZflMUW3eV3Yw0N
p/QUOPNYaDfGwV2e33zleTRW1wVCNqpfb52Eir+a0LAm0cUUX4WUa9/x73tJwoUXhcIeyXSJM6W+
xpC0OHCgktm7OsuS8brAacwCmYEBmgmznsdvNjlEoInWvHvlfk0wBgcUtSE49DywZpNLghra3Ez4
KS/5Sfk6P6/nUawJEfjsXFjvXm0oyHzWjqwZxBQv9wf3zSDHVU6JcB903h0i6rPh8aViri07HrOa
pKw8TcqXfC+qEdbyCZ9n/Vwep1mT6KMeTvKBp1pIb+XsnDW+idIrlAgVCtA8ASf9Dp7OY5iObyAV
WThyzT51WM7RgnBqEkVgYu1KpEP5JVdRtqJAfup5Vs3wc1XFnAj3SxnU+Ad/bNXD+OHvMJ08fdUI
B/U5Hnlt/M0I5Di4dZ7Ew3OfOWI1d8f0o0xEEmqzOsvus7FGH/43X/bpPffN1pq5CUlND02DItS8
aQtetZeMpzij3vK2A22lw9qdJc7mkIMsfXVwg/pc3JgpDpZHv4k1YBqKyj2Ep1nHfJIyGXS9hfh4
Fy7GYJF5rk/KbDW//oXYc8KceGvQmDdRhiEMmCmIufGA2JcIUynxNra2c7BO3R5/y10F5zjA+cBh
UX4MVcE+Lpn7iORcnwfGveESdPQINetBZw39I1pCJNtbdxPmXcSiZx52LKtkofVwaa6Zo1kd4yZz
zMytTj7XvPtJOoJ7uXZTR9l+OABAERKGZ+WjdmU8kr+7Tu351mBf6ldAJ121VTo3MZfJ8rVqw3k5
VvzXXcpLncC1XW8sPULaIAq8kPZemqm98sH6snG4abKz3VlrNZMx2lkIZmNQFWofwLhjUQKsIjPS
28DteEnG7bzrQK2mR7y7FtOKd/zJ2EO0mOPDXAcpp6oVgOSySuIi2MDmYxLzoq5dj3n2PPxk9PaB
lg7mOXErxgI3zXMcOGxAACyd7QsN0GdVaYtiqjlAr/kFv/rRc9eKgc5zqSaCly4fcAJXpVCd0jkY
eKC+N6kj0eorE1RPsI918mDhQZOoUiNvr9jn6yMcS5k6oS2bCz5NX5iM94EetL+B1bQ2DQVFfW2h
rlK4IvQZayiR+LWJpYqCkS62v4weL1+KhrpdT4AuTRS/7nx3xesVs78JLjZl6E4NOPeamG4Um9CV
/qZo2931/KnrLU+vP0H/K97AGRUSrmztRcruXRwvEzBZIvaeUlgpIj37+oCuNvYvoRMp7T0qTvkp
lItXRu1/p1wjxRspzh5gsrNMRqWmwB9kk6jun7CT+WxaoLfKo5pFa9W3rDruBtXjrZ1+4Y3YXCbn
4cHMS5BATgY/RNgopbO6M0zFD9aFrb717SVoqcXQx/xzrPym5zIeY7gxJl/J4+gsqwSc6IqEyS0t
Z0239qSniI0bQgRlidC5FfNQ5g9VvVHS+A/2DB2tymFJFr8MlF7BxPMFNlHA2AQVVfS5sdEnmrGY
TB1IFaajCrlpD8wKQVRRLmnmRAsK9hb3+g5e03VFuiGk96Fb+2VpAkBYTLVXTfUkCN+TZi0IC3Pc
EHheM8zu12m+zLFwzbe+JDl4gMx6gCHWAotWJkR9QwOEI+2L+0nYBHQxBIJ2ZjU1ReAvB/cuSyBR
3lyCAsLtfxKObTMvoT9iVhwrGTZp2ewkftxZxy7ieOlSa1vuSUFFNGy3oUmK8GH7TBtlmQjCq5ZT
DlaxgM1IK1R2xoaD2WzBUlA6TdvP9D1wbToibTvZtI8mLFkJb3ufJmpbWLKf/gLeklNTnp9UmX12
fWnUFobp7v4Wy8cn3SGvdSN/EAsOT3XycUEzpjUcXkI7s++4zCkfvAURRM2et3rkfDxOtPaVLJO4
rJSsnjYc0oW5bi4uYzvMhAIFiPgZvI+ebjK9/nMS0g3l15rdg+e7mlEcg1ylqlpIhjFHkXhIjFHs
+0CMUwIeuclInE5YJerrSN/2if9NOmYABT2unTII5gwqEsOVYV0YuubQrl3Yi+8E7HCqtkpYlyUn
AS8Dj50nO5jmwjbU7wkZNe6ldkfNwxqiXC6qGPO1BeK1Vw69xxBxDlzvsTZVhdzXIyOgMuICz+Pe
5AsyyZu9Xvcu0GpANmIQV/COs8tkdeMLkovM5gketFHip+6QMlasAmjDDhNWINSmkZHuivWUoy7h
4BGUwyfxf8wxAD7oj3VKSNnxbfIA1ZceOLhIdA+HUB4mgTRyrLOKZ/X2jTXSDk1IY7pSc/lWr276
MWNz4msQfaB9CWIe+yZ/+ha70a5cf3oBCCJqmzMRPQk7D2P2cmfs7FC92yC6GFXY1t8IgRXwo0Oz
s0ndPUoMw4/mRhAL55uUjd4JmCGg8gb8UnrF1MGtK6Cb9TT74V9o52/nEpMzJURPDJBV/s5v9NVm
+Hhj+93b81JVURnV6PsBoeTSsBkqDH0qrBJ+aZ+v/+pubxbX4mbzEWkwnJYVaFbqloi+ygM4r6cU
bzkLM7HiWbQEkrm0AAFsEcX6FudtmQ7J4tbGGM14jbfnzt5Ax7MM/BVdpiO9iVSKmbpmba+tt3GD
y98rAy/4oQwKpKhuVpCBoP7ARfmHcWO67ihKQSA+fWnr/ov6OQIh2o1WjhekSGrKqe19Sb7p+FUy
cQfPuyQlnsM7h5Di3zZJx4e1Swdl3d4saA28cEevF2r/q6P7I4jKWVliSFg9QJqaZnqILl01jM1x
uj7C3Ub1U1XSIWIS11iUXk+3UX/aglsw5Y5wZgKFkk7sMgeLLHyEh+dj7fnX0hf5cldcxbFg9+tD
+3WFtW9lO++7Bw2L1KpfIHiX3G4QkqjKvZttZVrOHge+34zdOUTN7uMbmFu/iu7hREdu6FNa7VmS
94T5dTUAqG+UUhDcc8kMAz9nb4GBFuSrgNFyDd9LNdXw267OXsSBALiUXP6EzRQP5mnoRRC7DiDu
ZiIs21Spnc8An7f+F7pF27K/ilohnADYfxqFnMHmOMiB0eKFexf17uhztVmCBHtSfI8VFck4EU1p
0QLbr6zqav7X4+SVnlnMGKRsfgLBi4GD8ZzeNFFE2yJXLV/H+oOrUVvO/7i8XQjvLsW7ZAj29Afg
FCg31R5yIqAoxiY+M89ESRBWuG2jQSCZEx945N7o00tXkaFuHRgkdCnWm12CUjio4oheQPNXJ/Kn
cdVudhTDemq2rHv0EaDT5KmLUK6SjhZKlkuLZFdgzkG2gcD9MDmZEZbHZ9WLmUxVV9OzoHtnm434
uuZlOWgVlW4X/VaKBVAzSLF0ZUd/C/GBDq1mbQXzUEPHRxNGlxorNU8gl3XiLLS2uGlUz9MpByd/
KXafnkTGUUy433CVT1hHB7JWs8FeqhTm592yFQrFzTGeRZXsxbEUInop14LhttSbHVDyZnKxN8cH
UiQ2BW+/EcSiwdEPMIgmeRD//EldR0BOOZwGWPc3lYqr6BrKRa6RhHjxJKmFtq/ZJdaR2UV6Eeqa
a7LIC9QOu5Pk2lllEwRyC7ieAw2JfWreHk2sZ2sDY1dBmhZe0G+ltEIyARy2NFUuiS3RbXT99GId
O+OETMMyqlc8rC2zDpVh+SZesmwcdClaHzwc6dUCIbMT/pRmuVM42Q9to0R1nqXqy0zyLuryUBaY
sOK95NV16501t8wC7+I9xeOxHrfsD4e0Z5b3EyHapG0ymTtNC+xHSatbVWdpiuoCHf8PtCohn88Q
3eEnWN+LG+Xz546Jcex1vPVHYnvkHBj1UgysIwnweIFf3AKBZq3Hli6X0WzjTShzLbsm9cpQN5zx
Uy/rHJuRV+0+kTRZisO32QBgpNizf0CKDK5t3+9itBnh+VldKJ1BHBabge9ZtKuey3zII3dw/jWZ
+hkX97034QATrwj20kIwYqBRg5Xqh+WNRtY2MUsjIhV7Mp00RBgtb9Kpf57klhBvfMk9WUqxebLH
Dwe67dE6cUue7LYo9FfsgNXzTYU6aJzEZsTUkb2J6XdM9h06f/D5nuTn+X0PU9LTfprtynXKp6EV
c5g/mSCnnfmVGI3tuwxO/zKqNPtmTFB+HwWbemNHTZPZKfZFwTkXsPa3ldUzS8kJF1vQqdkQpOKr
TltZGKlRPr2lZUEPJ+Ahg3xOJerw77cy2crFlEMzIg38ILC2u324nYqbC4KTKr99Gn6jzJFmIxc0
6mejWhK6eZzoAfk97H7yHhZxYf4RvmDUfI4GG+HQ8sZ3vYSmyxC1xiC+qfx3TGe2I5dPQXojQp5d
ZN+5qWqHFTfwers5XjmCUy1sk46VAPl0Uw9AqnVKX+VAceoX5MRFCrkXzTNYJCgXrqOjevPhLB49
Y0MeXOnnNdLVxmW02tcrJCpjp4ZMRTlYsWuoTPTOMyqPk8/nyRljLIzcmdhdtjZ0ZYMko4Kg9pxM
zghZyeTW5XQzFp+fpC2RqKLHAzRKS+89WHA/A09ncFdScBvLOhIuTAVajI7+yjbtzQ32hugAEm9S
FaPdp32+Md/ZtbNNrFTmEIgpla/ESaLU+SGs28hQm2rqa4HwKZeazR9YXOGdasZXe4OaWWtDBsys
Tn9pcdX0XHrwYvJa2vdDdduqrcHCJXAa4A12/7X79DajQYX8z0g3vmQ/kJqMYkFWSWtdVo/0cD9Q
cm94nLOBKME2NnHhjH4TFb5OC/ggI/35Lipcg0tcrSs8zcL+0sFRQg+GeCVGx7EK/wHZFqFjijfZ
jvYnIUr+3Bc6WLfsAK3iaD9AAopozJmiKlsx9UqIqzPev3zPle1S7Cc6TXAPMOVX8ZDxanuuavMF
idcpYT/lGeuFr2hvcWQHoyfs0WumL+GlxdOwX2vUxIMj7KkNhTHYnBRPtDTR0SdJRjJy4SMvjSmN
dOXXqDlCi8/hSZf4aphwWenCpnb9qrVpN4AyBc/GZF0q2iZkY4H4i2Ysq2sAlRMKXpNUtzS/mFdM
65chSErCSymBmF1jcR9YDPlFSJhQIeCMomGn2hG+HPC0t/sYIWAxrutcMFlcI/l1KGFLBSQEfPBi
cEm+aCb0TH2tMw+d5mq7sBqn4tf7Am15FebRNbPMwd8jl9MpBoPLqbN6m38UvPr1HniUlZxJoP9Z
JJ7+/x78amw2AQS/uxY8Q2WmhNiyCWOtr1nZBDPbamA1vG0r6XG2fUmM8DF3IZ5dHU84voUX471f
cAPW5Ueq6Cxi65E6GUpeQqhkJPOTfH7CIVmzMyX5FcHb0ia8C/QPsr/JcEchfwc4hPjQUIllonyS
RIUOgqbvtBL2ZMT5rNHXb73gGn7ZTHcw2npVFA06muJ97Jf5sUkrs2mmA5F5ICikDGdiJ+PHfTfK
z4PVIrS6cpAo2ZOB2a4lun4VISLODw8KH1II55i3Dxzww/GCz/sYo1KGF34UROswf97w5nzfgyG/
ua/fiqF1Uk2u9hPstaNjZ3Ny77Nresp8944AQEmbP/hLjvX9LcGH1sF30DGJvmkvdDIK3XzuZd+v
yayirjQkttCBFldxw6DgQ6uYvHmWDyBGF+dDJkOY/GOhm6LXYpSvTl8CEYRTAgs0OiUXbdEU8tIR
AMrk2TWino1dSMCv2kWiMI+wbILwExh0fRBLBicQbJwduFlBjqMBunUJbNkN53m6xP/PTYBQKEJJ
f3Rj6/ZI5/afevlkerrZiaizznZ2iWFso8SSdhwLacdiJviiW4KZFgvkpAjfVlBzP0v3+0wh2QWj
IPJqzN6lM+VxH2TW8UYs3RgOa3GaM9ap5D9CMN1Z4gWBgquneHqcJ4SXSW7YTaRJzSnTd4TbB0JN
sugdlAI+JZ7gSxKvILthaJguwXNydnFhwkOe966zNkzziH3XlJd4tO9YOkb2SkzL4FJK6zuFwSCx
HN9KG1pCr7kEs6GHk9g8+9phyj75Us0M6KAw85np0aA9mPk+QjWo0Ta3MwsbIiH7gG1UhBqIcBKc
Ryq7ccI4O5wEjmFxK3xeiWuSZ5ahQtdDhuO/VdO1WFKo13baZgtaUp0tcfKS0BKEY4MxER/ERER/
kQ85Did6f5hgy2ZyXA95bl5xwHtccRaYIEGx8JOPgjgYlQ5tXUjlS43B42u/asLCfXZcktwBGDq5
+5EFJYZQIMRlCdrRhFZrW0e5uBqFiarHNk4iLe0opVoCXEyjP58PT9eNAknzbgtsy+l7odTWJkll
mFSlXUoZPEc5q240pky6IOuvdYSZwcetm+HJZR8eaYqFov43aHncc2amdkQOIaPUc5KVp6WyCkQc
lGMysWG4aKAtAm/mAPV/t6yq6CC5EhIS1BE9WdIN/Sm0RrR2fZPs9ssJevqoz1YgsS00nR+eHccp
q6nkWMxbn4dB7syuc7lWDzWJCgx7/luxpYOu0gkQH4nGOf9jaEB0xtIa5IiBZ4uj+vnGi9lpCSQX
XIMQzxCylnTAvM+L5pc4nc5pM6u0ko7pAWB3JcFz3zrZRPGBCVzbhMl1o83BUgXSyUy2+pivLeN/
AwiMqpU08iVGVMMt9rEWilM/pBuxlykXBM7Xsg1KmipJbXESN91n5LlD9+dnsPG1IL3VtTJePGAz
PtN1khisC8wylYVfXbUKkq4U4uAm5YYoREFN4Sdy20rz4C8WmRJ81ADsIsoLYzLOIPlD93iv09gV
F0feuGg6ce5lNCuFoMUJXymAAsOJjbQPuzz983scehZF+hZA6Lfy8e+BXC956SBJV2AiKxN6BPXE
dRasmK/2X6DP0qwPBCk2oEGrOZiS5s35aeVNCLCpZVhohw7f9dknOfRKGYmUBtTu/vdrULUssyGs
w9RTMsuoGFm4W9A1NEtOrwntLekDSzrXlC/iR6Btk8zfwE1DfIyJrfX2mZRCg6ooTgLu3juY7w6u
vm9ghT/pbcj9kLSKvziCmnyjIiXKAvtIeMc1jj+mb/HmKAzgWeMOWWRw/iAnupVYjv5Dnd3JleYk
JSk8exumwmXSJpm+8ATH/kI20x5Km7WzqTCXCR+8OPbiaotZzNF26+KDHw2reHIwgDc8guxh1ALm
+p+NidGS3N5fzZ/I39XlnBHafRsbTVPuUdpMzp0/J0MdIYZHDRX0ig9ckDExxfTAAJqyj3TnBap+
6BEEo08zlMQRAy4TTLKD0t1P/E6kmaksnvSqQlClXooLAAGcKEpqxsIaVjjuDLMrZ1cxMNRiLTJ9
MzZkXqTw77JoyvXeQdfdNS2rpE2xhLEVaAzkj72nKxhR1BD8ESuai/PpxS5+aNRhE2CV2yRfLPv0
FVgPmpU1TOKA8GUNOQx6lc43FuSPyQE1KqsTXGvKmv2hCUHdgQYj7IvYPjiRzd/V2pwpJAGuo179
taKR+N69oTYCo8HnqvNChSm6SGlpy9nBplMp2kCXPUEV/1cfYDbqeh5N9mS+eBLR1HQ6ubon4vu7
QdUVO+XyOTHGxmYkA1CLb9yIF8IxVp7lmom2SY3kovX2DgjmXtl4YvbCifmO6JdgG+HA41ICkDM6
XCOzIoiv/oAXuszOujHf2hnGimfOreTAK1dYl34jEhQrdLAbB9u0puy9sIEWqmBO6KJ3Ydu+tKDS
KsN3vSRWeAZ7/9oAMFhrKOU9oUmf8ufpjpOIuefLDonnte8HsgBS1PvwyrquW9eqgvjb7N/5ayVX
tf0rwCfOUKGfa1698OfJ7JsXyMfolW+DUKUkR1psOodqgW12gc1YNMkEOLXqK3qlvkFvpPOXei/4
q1uWk+MBkPqe3Gp3LYB6am1037K2mBqhpfJZ7aVLmbt4C/jQDFx8Vx7yn+CrRVMx1TnGHF+xjToN
seflY5hyMp+P//bDaYuTYH09CZy+YjF1Vy9PtS9HbqiL6yGHyA27roko05eJMTLPsVUzCpHeI8Mx
Sl1+UxSI5cFyzBFhHk/4uJlgVaoGpJW/kJ1TGXpglQt9yVlNhdC1+kxV/FCGMTVYayDBE1usoIJR
DbGZk5JXUIGdiTOM2VPeVs0BCyamyFQ06UronrpKHo4FWeDIyZGJ1hvPiZ01UQtTkM0EtN74GA9E
Sq5SJPcKBpZ8ZJZOD8Ke8UTZus8XxwDq0Nf1Pi39YYXuy3urQ14R3JlzPoFWEL/ZtP3M64byRWJE
Ocq91uCp9TvvaKhcxC3NZ/IVTSTcfoeb4cmBPTrSdc1HXVfRhVCn6GRjOf26S1dqBHG25HZYuRO5
c+oP3HYPqAnYxtTxuFApfAs0062ULIg20xRPBM36AFgrlWHrKL3GxNWtcTXE503mAk3zR0LZ8ReE
qlBTWg42AiaUlJzyOmFSGTGJ6eyw02WSQ39HlNj5Q8OyTEp+ynymQaretVyjtYkXe/DFXfcHqIVV
FSAcFqF0VeIU+0oIMgVqwN5/X3TVI33C9oILkPnkFUux2kODA3wi5v5phyej2ysBZgkhCXSH+oof
N0eWaiAaG6uNmAQ1TeelAmP5pb8tjGKBO4A8oL6Euv4TlTNZi1/Z4jBpeZ3FSX//TnmV97F0fN1k
7SIYLOGN32KyKUmqPin/3AUriyY0yTKHytkZnarnhGOQTTK0B/a3dppT1mMmjz+LOCAEfOm4RW1x
mA3H0Drpzh7ybnTdvC7468ce9ra0SJigOXmO9tUj5vqjn1/gJk7pT5F0IoOEMKO0IEbBYpe+3LuP
BJY0AuRXLzjZmAujCS06LNmZkffOTAUQDz2j5ZmvBpUGgnfLX+5+fUsrC9s1wSIzEf05gRZjmF0J
O5cyznKrSTYbGvAayEE0B7q1RnqS8hrrfm2u3/u1wFEqGvpSbqDgo3zep8KxlHzcGsDJrgyNXJKu
9yeAdzr2PBs9MIcG5ySQkvP+7HcEYUhww3Qu4nyA/q8eGzGjNmDPTOqH+LeZNTkJfn0h2IWgKGUw
eUh8bsxAm6+38TEjfIR8IyyDlJKr5EkoSZbETImM7FHiU1XiimY5luxfzmmQzfGLU5LyIZooA06W
RXioqMFldRfrDTKXdmKcYrvMQIdybk1C7nPZoyNl6ZxGd7dB7Kg5Y5JZTRz7U4/Nswff55lhSXYQ
WLx5DDCAXlKry8ekOpyWvHbDJ6LB0WfhXvh7wagbhgl4vSJcDGfLNfgMPzqQMMOnuuXIUlRhKKzj
PlXFLU2IHeIbGbijgXVwCC1rd14y3AasyX4CMkyoyNIk95vkp9mJupGnJrVsTmZS1zfs3wTvunuW
u7x7DjqWYthDevZOlKCziXtxJZfdpxW9ZX+TO1ITRCB9Y2QEuAOLluCtmCUJAocR57uE6/Xsfwoo
Ws7IpRsbmT3vtxR3OmaxLy9f5fJ3bTxNx3EEe9NW9zoV6ZWwTU7VegfZMEMgR3ZWoKD7frF/lnJf
lOoLiP3IlAeU7isokYCYLeTETjKZtU/AEx/60cQ+0XJSqg6i7uDHUqlEdZ8epIk8+VZAFVtZMZAr
Ct/DcJYgKWY3FylQWzsB2+czksAGNyhfMeGp8bkKm9tXiXy2R0nJeN/9YoEVH+ImsGlWJGuuSzqQ
91KvINIKNqZrmqGvXjKMXL6mWKOHGX5vYhLOM9V6lqVyO9EfRXvnvCw5bMgSGZP5dJgAE4G5HJ7C
ybNv75otFp8BLSHTG3pbllZOmCAdja1LpzHdl7QD52+z/Ut3AfZiNk7veehn4IGmfRozEL/V8/iQ
ebhF/vPoSYYBjdsdlRS6UEXnSzU970zKv8mEOaLbwtk1Ew8Pn5RZoBsOvG39
`protect end_protected
