`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dha/a+q3FYn0HVlark/dL9eKG5WFTs7ZZirNn2JiZyMDhD+yVf6YOVbeSUTbB59BHRuMRTe4HzMF
fb0dReVcmA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L/ZWUhD7C1wMz9cuwn0TiUsK2zqZcBb7ft0zqxgdS/DBrX8d4UvO11L6mj4hlqYr4eSJsYayZYx6
9z3WLZv8ts+V58d5ow1lZp3/rBgg5wjNmEtVwPtkT36Il0TXjKVXRTRW8pgujZHbRCJmMdsI6ehy
B8jk5KaPa8BeDG31V90=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
prNGuml44BHYeOlEWt4UF/G5iqeBKYcKR7cDC7BlYe/+VQgAgOwzFUiQuH5qGN5IDtkYAw8fUWsX
DBY/QktpuaiTarC8x1H8FtTW8djc/WMz83EefgzjSPC4CfBmdsKhajVNRwaIxkbDn/m7DkNIxNqg
oGsIhNJM64YlEzAjdlsKmVZGh+C8AeyQYt3R6xKX9VX8phgCCfKWd/6ANwOk9zbI09xjsSWAlSny
KHmRF7eW37kBaGZmCKX3xWvo9ysIyr00HTEmf70GRSVAwdoXTdNM18UfxDoNNFbRSJxaAfmrysCV
B0L1uPFmvdZ0qyInVQ6pJogDdEyFJOWOjw1D6w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EUhMVj01KRu+/d1BBnp5fozTKNc/iLzWR4cuQvtIjp1S4QppFBQLbv2niR66OIEPXGtWmg/C3bt7
S7eCJuk9ASctS5KkEOkqBlpP8QAFxBKF2uuG498unR+eG/low1R870bxI4+UL34+zpr1EBzeg1D1
Nfge4873tH8ERTI3EvM74yfhDWXR920MVAjCjBFGhJZSPrmaezLuvU0R8J2SCDMZ6Pw8leenxQI0
TuREcLnyLoDq1zXvjKwzemjPOnOH8E1CnfSKTqSyDLB+JZxvrMRqbCqCM13onR3UToK8s0Ii/geI
hFZZrV19JyfFvi2ZgRQtphySmAkrVv7oC29Nbg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SZFp62A/hKMXaqF+tV4TShGLMAi9E10qKJGW90/3jo/vBfLg7J2/TygMjEYRRy7JvszNgUFzY3LB
jP1rRKBpyan373Hbji7JayH9qj12Hz42uHNRQV8lKi1fHx3dsUU6ECqf2EHZJESSgAPeRv1gwlPv
mV/im1bLSuck+d21kO6pljVOJ0J7IAgNyx0q1pYq1Y0VKvA7sDwUAXPdqzZj6V8jKr7a1E5g8sgc
mgDBJzl4deilCuofpwA9fOKlAG86EHAm0QAZ0XAfih1UeZWn69s0y9vh4bBCAbY7OAqOpNfVao4G
FrcEywehMzx/b5V4ZXvUi0zO8Y5UjAXjbv9zYA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z2Bx0VTdG7Pi70pLCZP9uAOpM6jUBUJp3Ta1oJGurka+ma7qif/qxau8roqJBQtxRrM27OzMaE97
B4rcIrDF4U8IePphJsK37PQP0Yz2FByrdB32rjTDCj/2VpN7y1Z00JZi/35AAEn6fo10PlQ60zgT
24EzNmwwUQ3P7cQprtA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
feyINVT3xMfhjYK2dAdC1z/oYf/Ff2LPnheBDSSHmA5HbOuaEPmaVBN5H07klhyn9WUoSOMBoVZ/
wESscqFjNF8w7QIzSLEqvFj4k5dMi+/iV7e+Y/xsWW+IBVeuluuoj/N46erURJ7mVNjalWHVYSKN
51nYUOTEw4yuinyTGpEMM4X0Czvn/dMd1xi08MnAGAk55o97PNlCV0359gXOFsCEqKlM2QMp4IVP
qfOJHW/2oOOT4rVUMeTZ8+S7pin7ngkIGY4QWMfVl28l32xd9htKk4+6Hpc3zopZabnOByA5qj8E
02oLYpWgSyeUzLnyLwrCLtyuAYVn1Uiy4+XvKw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 308208)
`protect data_block
xL0fux1EY00x74Eghns/k83ZBsT9T6in3BgnO6HgGC7bRIqc39gdiO7MnKLk5fldUQzltLOzSTp7
RoShjiP6Q+gxQ+alOQplbwLAYs/bKL6bQz7ELi1avqlCqoOp2ljf6dER23PQL+1kS+ss1iArEu0l
F5Fabb/d7HaqlXaXAgubC8SkgtwpukNmfwbx1QlpVfOFjWZM+RiQ48Boi3ENcmr+tSFMSXFPBSeI
IYIaA5nl2eiwmya/rLlSTzBIMQOzfOwuuPI2XKIP5B1253Jg1qQM5oQ6F9sUanwMwmtE0A8bZRBv
slH2sNy64Yyn/8ejrLU2mqYAJYQtLE6BW7/KzVUl5Z2Wr1SrHccsOixk/uowoAjONht+aNYTaVuM
R3jIjByNePwC3mnfhjouxoqW+NezMGoTZEktOmVAb7cy3jm+2O8Xq1qJw20FPiBGIFsqYrr5oaLG
vwfiw8ChYK+vAYvaOLKn7++1zlYdbpeUkCEM3IpfPs7SGLQlRQ2K64UzZyVmwnLX47RciQQon8li
nSWSVLhOzpInusRuH2zaDykFaT1fsByvVWreRqIk3vIyqDnmp9K21SMcLaahgf3jNFt6jX3INCJR
FpVWAM8ixfyAH9ZVTPBs5UuOHbnc5pIPXq4VvpAVppmlFCzhpCPg7C5jNGrlBT3OfYyiPO2GHokK
DjhaU2rD/4Yb3NdIDJMHYrUF/lk3CKl1GyqNLoZWmznYN508FNx4P2Qlc9nAp1155PPE8vG/5gsL
CVdeLiPhJRlblHpa87wClsbWg5Gt6xRHk7M9UByxA2neyybcTrvGWJk/+RdgYFLvVPf2WI71Hmo9
fKS++buX0gT51xVR/Q+AOvzSnOu+eoY8L62HY41ZQsMCK+mqIpL1479KzAdM00MMFC/V5nSzg6Bf
KsfUEaFqdfBZUyChcBbvDrsOcMVUHU/JM2KSBbjhwMpk/LpUSoJdw46V5/eGyza3deTV8kp24GKP
x8NyWv5hPhiPcjwNqQyo4ZAStAMW3RBmWtvwZEmFp6tM+h5h0lhnyOOUrlCb2jfrq+JzNdzITkAf
1j7YrULGLxQTeAijE+tLsPGDVCbeJ0yVBlYFl7yQCoUt8T4flbLg8aZzi4N083NSJ0kupt8PKnFA
Bm9vGI6aKEBUFqorK0qrvfxbGgzoEIY/hqoPov19kEl8cx/z35UFws6l+o2O/JyobBAWTU2FSjq5
GbWzts2cDOlKmjv+LUR/Fn7vlmm3iWMvXAWAuYf9OuFhrDXB/8+rzLhJAbHfOxRLublxCU0NwPXy
tng7as3+a7B3VWq48PlXdKy822yli1HNYjtdtaxw/LCvxbR29MZ7tSsHK9NCwbz4e4HQALQrykYB
809zOWQoW40/fGO1fK4DR37OJaQfS+N3YuFF5xG/n5ZUbXixddzs1Vitc9/AxI3/OMCMpYNUgCfo
guzO07TcsSbZ6+yEn79qSQV3A0YkVBHHDa5hzsqTFB8EyCRggFsiUJjT9rMtywS0z5P10Wm3pTFR
F7OIC8/IN+/jSn7Vfd9tfOHzWSyO0Odai4cU5plCHjyc1/99/UvwHLPwDNOrRIrYX7DrZoTWH7Ze
DOImf0mN87X2Y1qKJGq38c6Sg49xlTH/hhWMPYg502TvXiqFKHbFXU50+cO8QavG+CmUdg0spQAl
gzIZPzpELU4dWWA8x51/EiwNFoukLlOomavjDTWoGaBMBvPjwMM/pHOsPCOJ2YBCk3eIvvLC7hIY
vqGyvlZXzNayjR6cP9VSyT0KvUGidg4tHiNljzkSIO3lfzqNaudpdYxs8Enw1c0mdB5Mch8R6sMy
9bfW+qN+jHVP7e0KO7Ts4XbBK7cLztFZG8hvItubYB7q/0GcL4WiovMDLwIncwDgk1HfxYcOiBXP
c4gohfuuagP8FQrYiOshY96qCPIz+yCCLmwX9L7pkCqrKI0TPnddo97SIjKzMi7Ycqu1NDBaXbil
Q4kuzA0OHSl9EWlde7YZHevo1Hzux98t9ltsJ6thNiYPM/piLGCJycUibsgBgoSrrTU9rypapzL2
O5xYt6h4KU7p6cP/43bAJTjv8uXZWk89FwWz3MprXKFMuCcZhQmZZfIJ0sAmKAD1Qlj4o+yL6yYm
d8Qf5Le9Y0rhdl4QfK2WBBqydpIdTrHVCWDaeWS3X+TIYZsm+YrrEwv0qZFrzUzF2aTr2aNiS+ZH
oEgb/v3SioY/CUoi6xdpWfHGvdWudqeUMi6qYBVfJMDg0tmqyiy7M3pIhuezfUuFZ/iUBk1ORd4c
EMbD+k4dO+qkx+/UwfhRA/fwTuwdwy8StF2MxO2/jysz9scD7q0+IzH3iBMUSvMDMvg334BZvLQH
a0+ucAV9soMkAXOxkLm5H6p3EiKJiIIHM9OtBpmVKZ22GR/LW2sxE+uWKGUd4pJp0DX9KKjX+lWG
orjPp4NuN6g+3qT79g5ivuJMyEWohvkHke7tgE8SyIauc4hBeHvOSb7igaUf8eCU1g0c+6NkQza6
qygsnW6P86JFYEx2NvIXi304mUGjD0FgAVmv7Yc1cEdcEiTTIlSOHdgl5tULrbfnEfIl3XfaBPW1
+8oUXs/vfzFeh6GzdORHviSI2xw/dWwgbks8i13pP3WjpntP2MpoCVoveXOrvmnck/0Yby/gQHkd
mMevqY/o8ED+FraPozr6Q9YOar8G+O7gZWSYzOibwvKQ46o2PKp4GXJ1Phg9ziUk5HwYxGq+/uAt
l5X3f3Wa2Rp1sC2Zq9RYWJLU2RTP8OXH1T23v+2PUzJjhzkir9H8VN9pTNyYd2j77fcNKtVOXyZi
usw3imjfRSnOoXPKBpYiylFgY2BYgXcsi1Y4UazV0JYgnm+ct2U06cwNOuCFNLgXxjGMgMVsxY7B
aKvAKfyO19uWKkkC75pE4SV1IMKqhw8PxueEs5A0c8i/X9FwU1WG4g1BNpdDKe42OZef6JQxgdgd
dhrtxjNQW9P5+9yc9ktRu3yHgxkOo/SKWtl2VPD+Cp4670Q4aUu2bKS1nBMwlO90apblvVui74MU
/7p4DNEbkKdAwdj80FFOkSj3jHL1uA0OiZEQsaP9UWzM+8U2uPr5PdRh4klsesOwm6prcY5czlN/
1SwXFa448/hyOkAsBZ82GTtJqsbTbOHh+GoFt88ymKUKFhXkfrUsaCvcQkj8k1U/OTal+XnQnEUT
odOF5Y3BUbVMDOdme0mBbxHzY1Gy99iVxe2S+JzSnpQT63DIjUOkQkfbvRY7CVy36HMTpqSiC3im
j7SN2ovv87zhvVuJdaWINeF6+lf73al84A/TE9Fsd/+1rS/c7uBpqnwpJaAu+IbbLz0Mfqp9osQ2
h/lKGMST/lEz8Bd7SuEmJvnbUXTmrmIInewy/hgVdvkOGhWT458GAzL5KEg1O2WYKKdbfucucGYD
aN7u66tCV4UDskFqdEuEMk/HJwX4yx/yhZcbYzsnjxV7eBhmUbY9gotnUc1ILz5xbIqsRhFlyZJF
53DCpToD5sWq+T8YEi98KdY8Vv2Pcpjyk3TkBokAQFIKQ6acekPbdVMIwqVf1MUA1eaEyJaLhrJI
bNkRdg2haq0bsh0E5efoCMkpoMSB3DInv+10Jw44KFqobqYdZ4s71p0OE+xtNok8YKNofYoRLTgP
GSvCjOiE7Zbz6+z9/9bEsuXxB2EYOFxiyiX5yvTf2yqkGm195+N96Wa6ienTxFy7fvi7ZBXHG/UF
SmquVNKgTPpoz6CByrbzEPA2laQ9cgYadqEPoHt8hS+iL559BaoTmCR5VCO2JkSa8+r7VpKMJt9x
Dlx9qHQAnpQTOSBEMf9/5XzllVFI1H/vqMEKIuo0R4wTKwp67MUlWabNMblp7gYn/6KGqaK604tG
LC6fQ/+fK+5yTfpvbDpXqyoZArEYBO7MAcN/Fl2iNWyu880Sv++1Vf4HE6gYctGhCtZWZKQnB8XY
zPz3THsb8lCFo6K2ywADS4ra49rmyP0sABdn+GfZV/6Oqm/nccqFoVjYH5zEJ8dOZwV12MJMf8/x
0m7/Vn8ZNMBpIR3QhEtqQDvvZ180Fp4pB/s8K0s/xbM+VpGZMG6/tdcwQ/jd4N8rv8M3EgtkZDz4
Bn0kMRJ8LGTsPlZo07HKDwvRCCiQlmBAVEWMN+HuMhJjBJla93Ob9oY6liEb8Xgj66Szn/oTxEC0
YoPMD2u2JHboXb02GpX6FdD5sLBfYknRC1j312r/LYmrIBgqlbcuEwD0A655NQcJFvX7A4QbIKrR
YjkrpzwJ46gutiv+6L+zZxp0+eKVlLQ081SC2H9XtyQBA1TAwB0zI2er9ffBXD9mdHUZiRKGGScI
rsorSgtYVVDtpRTScEZbNQzoV3D6ZOUv7ubU0xAJoqe9OAPA8Yf7r9aSM4JTaH6IQwGLLU7j1guF
KcSnp/YZu/kkfme6huR3fUQLL+k/CNv2Vuaao8ko8erdF1pyOzJHhWhTw1NIogNnJHLbS56wrx/4
VvhJpQ45ABFcBZEsWWHM3AxFM2YFGhpTZ1aMHPyenIaDnh3UBxrbbqGzor5gu+ivxBARbPFAwEj0
M9Fhylx02zdefYyps33/MC5ylWE39MMg0Npe5ZXSlOUNABBEeGP9FG1lnrq2eG8Hw94UpPbtCt46
oi6V3S3IdCc4YvQPrvniATV/j90YhJrn3DmiVaj15O/f/lQ5Ko75gHJOGwCNU6h6tuNWijPMTB+R
IJ3aaC3rn1yIkmgP/MUVq7/y6E5MtotZIosHuCv6qBvaEd7dqISrlpCzlDf/jrMUogYnQb1cJQ5X
fc62Uyzcxb86rSPFy1/ljBkf7Ar408oq3fBcrsQifSeNfo1ciIAkH98K32jUGPhpbmHRnw1NQkrn
frlD5HlmBH+epNUwC+LhpO4zzsBs9v3pd3/s/UdqQ1gzP3jK9JbrerFzZ7hHSFKzy/KAM73BnQdN
IPBZq6Df5rQkAYlvXPIPRGXGFLKac4UWuXkWY40ddBBhrv7FoXL6g2YTO9gUp05TZrSAeK6SD50E
M6E8SJZojbizg3n4rI22VMgzR63mIo5GGrRc5l21r+bhdxSx3dqORUX+a/TNK5WjGeb88x53vdyW
bLWtgO5LgnETNXfXMMbDkB1pl3Xn2Ci8c4lHIoCxaSmFzQVKmDpGoNAlZyrIfqOkHOmB1/zPxgce
a5vLtnHWtmZB33EHQIrWv/7xUitbkiL9X8aEIMpeFAEu+xTzP4XliQHhUX8SCnp7FmOOK9Nu+A//
SqNwPHGuJIJTNpMwkdJh4feuPaquwgr8ouVr83uS8Zu+BBNgOd5i713erK8t2QSxDZCSLHV7hQYY
mvBBZR+5syUk27ZLYSO3xer3R2vLr/Bjl9pDJGDyWCS22ry5641+/fZzRaU9Dj6lhZueQ16IuptH
AkK+USOr7R9soRyAqbUG/6Wz9EZZcdsqbjfMQH1tc1+gVYp117Cz/OVOw2cJlTGAYyGoCVG1wRJD
wfDSOyDVdkVBqhN7UX2Go+iusjuJEGHt7OXjiZsMl6/5WMXaQMePuRqfdfi4i+VM7ScX/MvzjaaE
pKu7e+eu4YXI/RviPIdW+ExEBk415dz+BbHEtXwKWySG0ENNMzxHupJDutZ3JCqv53iYdJXCCMPH
edeR/xX85ifR4ui3vSH172UCnJT/VJ5zhZ9H6AMsh7W5T33LOFrae8zqklPZYcVOcJJNPN6qcRWd
dM8Z0uYG+je2VQuatTY/8FB22lWwqCYmZgyr5S/SgKcL6yiWD5o1ZtMcHvNPEShisD4y2D5OU6Ag
BjYOY4/VfUzfclP/13bV/LDyS8xrlilXB0ZTlb18q0fhKnXcatYs4yHSyk3EBTYSq7/VOoA/ibJy
swIssvwMHeyT4mzIpW/5TGpGsde6MfB1dk3zBqqmpmhNFovt2blbuztPMoCfNiUEMv4muL+tJT4a
CsgpD+75cafdafC6kzpP9JPhMcmXWxGaH8teTLOERhogGLJhXrWDoc7KpbnVYqf/pW3HTPueD3Y7
Q/w/0hNx35VmaZH/zN864Agr8QvMfApmJIRRlKAVC8eFzOqUad77MoJuy6Dyubgia4521HC1LX9q
Bw+Lzq3XD/C+MiVDb93ZTpv91I4K8YChrRaNe+ZUJeO4l5ghYtV62vofNnPmRSySHltqBN3GkoxX
aIb27Jx8EZsi0FuDypB1jCxakk8am870Fc7LXuysugscWhFIPhOv3nU6k7JfOphFhKwh/1ucF5NL
8x9X1aIjzZNDt1fAF0nv/jrOYUmRMnalOyfY3wS+4rWhrMuLBDffMuxsP2ux9wcch7bsC9+hdZ52
7h06eXxp8alPJRffsKannEVQ0akqXPE8XzvRdeS4xALl62NU27ulb98HmdtB5qUEJcHuph/fQU+o
ealWZrHpVOSTO6gi4rF/SMohc6yPkaFJeR/GRrjFhqFRRU+7EMEV8ajcszrp46cSmrh2h29oUGnn
0IqGc/WRvX5iz4qRn5aN63TfWajzF0L7Pb3Sxi0sJ83PMWRn61X+M86Tq8oRQlb7ze59597VranQ
4l657XXm9KJ5A4Sy9DZ17POyYIYiWXt/Kk3WD9de1ZMLdmza3xiaJxntWMQ5u+DSTCLkHdJMn3xE
PV3aSJcuUU0+Dh6X7HX5tAzY5Cd9GNWxrUYA9AMJtC+vPiOeCYCS/0P6wgVvS5k0NKc90EcrDn3j
DZBuaZ9XpoJHU+9VQqOlcYbU9oqL7uihS/tufffdbytgai72+dulsSFMK+jP4GQw/VIHAiEbhWjY
yr9ZgCbYzkVvNp15Qm0en8kD01qHTpTvQY12OgqWCFazdOEBniqVXuIlSNpKWMrK6rSXtBR0x0k9
CihChSBi50JoJtyMtzAH92a+l6bPEXWnXilkDn6RzCLS7brSSMukDFkZdPi7hAwn3NKjlDKNTzB0
yiK657y5DBraxn6M3dsFQ9SAYOygskkeLduDTiBg5C/ReXdQ/f1VXiM6Hrtn/RsjVP/lZe3209DW
NBs/7PdPkn2GVGP1r34zf+BncIfNKjIZDpzhwMjZ+JbfirAfPhcikiBdQ8grbPwMU7GYNDbxqDbO
9qKVgRaCbr8BlNI7UxxATflGrd2hL9F2tuwQCCybr2fBs0AqR+Zhmti4sbM/W3W/nsmrEPnDEFej
V0I1VahAybfsqCOzsRNh0FMRmGyVk/WZAlBJDrIvltYIE06l2NLRyqOAHglfVbYZJS36Yq16peO2
lerA1u4lNDWxbdGhTXpkHWY2fbg0U4PiKV2jzX9VLSM+uHHIi4jQ4LFQr+yeEZPu8JgcamVgrnF5
v7i/tMYMu2qkpXMfJ6comjv6X6MOZUELFwjjRil6ZonlyrJr4PcGr8m9VFdWwrGjBV+0hwUSjm64
VajXO/sEkn1gFT8a5CrQFcuM2VnrvEYVarPdkC1ozQrQ8Bfk+hmrv+1cdL+bWBtmuBp8MwpfP6qR
HsYRNfmnM2Cdj+xaZZPXKkxn301b0ZTIzxuEWqtpeOZzzEwZvjvscEm1Hj+ba7euJOCnM21/f1n+
SWx/zDi46JU8FcaTXBiF+TIESdkr20Ol+4Suo5bU1SAeVur9GIzzgFbiDlymRhzU9hIpzYjsrdCJ
9aiMrXCHtxFvhOte7vaKpcMM72KvvTnS00Jjo0j/NxqNfzOxJCayIQwUrdot1hHxUbJTWfzcconm
zGgyAkXTRwKCVdkZvPnH7mrBkwMLB6DtSKKz5FCph/s/d4uup7rQjsJv+YqvcatRtmIqHoYF3z5a
HVTeJrmZE1jdoszG0Amr9UjR8BX14jtT5PBOYSFgk7cKBILOCO3xVSbyEE4QoAEB1GeFkB4C1JkD
AbX5tzVk4XgsrBzef9/GiHI/rPrlQzXLU/rb1utVnq5/3fooXGdukmAOHVFPKJWh8t8P83u+qbGm
63IweI5sdUBFYgaWTVJw74NUdWbwv8BWHrF8BbGbM/acA43YKIT5rWf0o+vm6zRTaj3NGVMfg3vl
j1KrxxXxbbdgUDZJ31Q65MJCKhpeJjOmb9Rb0Yre98fuxYApr/Bw4bHOg8Lwu8acR+hXDQNQffkk
fnA5C/J1m8xP7ozlk5HfeUdEMgePj9BZUf4AyUln7q9cF+ydcoCMocCAPyAg2FOq7bELYlfre4yD
E9Cwc7918HBhKwb4wFWT4Kohx0G1S//mPK7n51x7yk6MRKk0UMB5rBtjlmAQeNvDNi6dF6RjsZUH
CWnTS53VEVM/JbxiYzIbuHJMC+0jfpwB95HmtVRlwhlhTgfweQAmujYOgXgF9ChGm6AyH4q5z/rE
rwboi5hbddFAkzcsjttZVdCtOkuyNCt+XnsKA9F35QCfrKWMTdRNTc3G2v8czW/v6S7F+oi4+8if
DNfiyHyHNWyIfkbVwweJkRuyje1a/lTLlpTe3fQ50x1UTaLz/tNpDz0GpmAZ/G5KTV7rPjnt+Wvd
yk9jal63BiAOs5uMFPlXSIlynEBk+tBQzCD0WgeoB3Ybn9GzPkg8DJTxjxCLlWce93pTRd58pUkJ
/aKLNfk8dj7GhDUBHBmHRbGWuxH5ujpo0RW4Kk7jtsJ/5Ambfu8w/X1ibecCd/8yO+xqB5KUv9c5
//u1sjulpcYGhb33h/zCma87fs3FgWSTHcUXMpkZQrEpd4wXzrJcgthy1H5U1Wrmzdxh8MsnlaQH
0ewIwmVF5xMNyQGBkoM9mVnDVQhUp9ukuWviGItpMRTneA/IB25oGz1CEh6vh8w+O8NM7ABvhWrK
LfReUnjD+rtmZt/v7bKxhVA/HqLAx8Qm7Fr5sk4lfGZSfMuIqy97if3ij+/ORq65eGY6c/56FLW/
Ru70ibZZLYJPYDMevUz4b+6n1KGFJjRmjCI3XnheTGqzlamB71bxLhTNXTiso73Rs2fKQiuxEikY
ZmkWzM/Ac/DerQVIL87eNmUHFI2Q54Alw21LdBXIqt+5sCJa3k4fKWZPwfne9AyzylDYYL/0aa/X
4JFTPLGbeKan+RhsnnL7qnMR+jmpqb2zNzSISpM/Dd1rmIvwCwQ2AE3JlEdrge+75SiTJs96nW6P
F3Gjd0b5NwBrbAYIj8GUrrSH7eEeXfVd5XKibUpagysf/PFFVJ6+XZMmDv4uB0SPjMYI0x3vRC64
/PFixMAjke+ItdSoNADMLq+0kVdrLwBMk2jebPI3rIHS8Zr7qBCivPVt+mzhoHTsTrWDTbeSmPPA
XVp83GBHSmv1mBcAdOIkG6nkxHG/cxyxutApOcztokm54lpjsSNVHgn3vTE8IToUzeKrXmXvjt4H
49VUv5VhJZgftIa6JrXSQ6jBtNyzAp0L5Gr5LW8EyQTFq9xPZkNhl7Z1eAVA9JuPnjiPFlXk/79/
n5taU9K2dF4SGbcXRvKDA/SKJk+aT2I5MxG2oNgDLbPS2NU90G3A/1ACxUrTJnL1wA3xN5EmIEaL
S7m+YaioowdmoYwXhxPsCg7FSbssHW32IwE4AhA8VlAP8d0+YqSMlaH/tUoaQIPCdWEkQEuqMA0U
onoD6UEacWWVjmNk9fiaK4TUxrlD8+eTRv8opB9LgjP/gUVf9HfBG01IZci58nyXK7jIFl6pXzRF
VAbQcmJIkac5Kml2RcTiswqgxcB30Dk4VeZ88AaMaLPzS9CXmLlcRM7K1QoNAyuETANicK5KTqac
bw4gcCSf7O9YOL/Qaxnl6Vge3Yt+UQ2J7rg1bjQQZwcD/iAssPGDQ2/Ixuv5Cx29t0kA57EO564f
0Q7AUbEDEcQtbHxjfhmArg2uXPEvn9lyofy8vW2yQQhMuVNN+IqJ+1v/N76M3niAe7nvYBfMk7Rz
jQcgLw+YzZCrS83C38YZ80Q3LW9kSl9RD3HZ9FjVFK4G3vQzaRSzrpjRJvxlhCJhLob0mJ0gaO/f
d7QFnKfBzHGwUsDOy58CYMcacigNgTpLhFjQIcPGx8F41VXqrfMsxspMM2lyVfVzP5epbC7tdf87
Ppd2Ls1hB5tx11mWT5D/flS+jk2moHvE4Qg35EvvlCUPcFQiYvSJAoz/BHIRN8oixfCO2AHQRgvp
ADjXCoho8yfvRL32DJwjZy/Abn7gLokvuUXIr6MFyhdTw0CgT2qYq4UuimQAW9lZP3e2NSdQnyfq
FsEZ9VJ5FfIkyiPf2d65dLy/FCxEgS3rq0qJG6NBiDNQXBNgn3lPsUlo5MQRbB72ai0s324zOICO
+YcMm1DRwVW0bYOIH6IsoYZZjtMVTKvMlAPnECCqEa0LCeAU9E7EXF//qkTHL4G7OxVlILNSN5u3
zLVpm638AcYZNZeKbd0QxKISgrCazCY1NrMFkdxG6ryUo2pOy7QSy+EZQ8m0kAscuV6K/TMUgD1u
nM/tjXXEMw+aby2N1aEiOVohXvv2KNIfkvam0mq8FLsy10J5CAXnwfX2FP0E+G99q4Ga2t4YdL1X
T3sup8yBX1C1cXZTuZmxPvLX/p7p5j85uP+bf5cKPfNqw9beOUYJG35CNLBf653LWVleJbxnH/mV
gAhsXqIWcQ+CTVxKvm8iFZvIf+UUmsaAnTqH26pSLzKGJeE84BtdNymn4tU1nekSzJ51C/xynsNk
0iYqrg52pF0hG2BUk537B6xMtbcep3HgIXv+u5HwVp5ikP48vCv7bzm/VuqV8KxJeMtZInB3vP+9
Vwr1EmV8yzumxWuQnfkEbeMWGApl9BcwMuPP6bKkT7jtyOfu169GuAaMYbTSJaSzuP2/6wOxl2q0
Cd39b+GiRXzdhkK4SVMjwr89Fy0GU3ujHWsk5lKMxNSkR1UFdCt7FZEHsu3ESQAfj6xQoPUyNl0T
WuWpfto76+2lkozgw+q1oRpmsayTLwZRL11nbl+Yqn8KWEYC87gGwJiVLFSrSedYj6/bLVfBlwKj
9ob+R4iMfja4nXO0r+izlOmtr3P4iz+n96+L6obCRrh7nuiEQpunLNDQRGmVNf3IvOjA3ybAylTO
ZG7ool0dLFM8HV89+5Tw7n6y6nw2JCl2ajvl0H2ftCMBUViN4c+puCO1VLR0CJv5AfJdHCTWyXsP
LDGlgLLUcSrhOdqTpAb3kS91P3MhCOOi+Tk/NVDJTlntxfcE+vIVDoGycZlAksqyqW8tf1W20Q3E
wCSnvACCns9voYZEyGSZkKdJmOJ//NU9TA+imoSO1JB7NI5Fo+wSNNGUC1PmHriwGAYVvC+J0Ig4
as9JOp7UPAwk58H9sj3c0D4N/xF4HgPqm/BB8jzktrwKJIKQbfS86pJ72iOwwdJHY/LsyrMvkMlH
VqnVBq4nnhfvytuiirNnMmVSqXNkg1Ch9eeReA0InxNcdR7twWw7uF8PFpk6tQD+2E8DFKMPo+AR
sOopfGHtKpwjDUwDcbIIqv717d0HRUyxVcWuaW/XE7W/nXZjs9HGIXtf7CI+QWosiqQbgl5vmjli
e0bm5CnyePhgEO9tma+6XHqaVGQBCde1DjCdhyi91a2w2TNWbLvUB5G06ZJ85zSkAnfqXZHZiv/E
F1VduROV/mjD0d0hTJLV7w87YZoAkNpjRLRX8vFeSOQfhxi9IHtljklxAnfPFiPNwC4lXuAqCItU
MfW96J8cXEzxt4yMe3Le83cwqk+Jt/5H+fzNqHdrbOau0TQNZWpLwww3qdwblGvYyBYVR3xgbr9M
C7jo3CgSS14hK9FGjahhAfgll/Q19gsdpTz9z/aHOwZV/bg8zYqE9Iqg19Q6HUlSs5c5iDyb9j/Q
q2e1YVBQjTe/D7QhYjKaDWI18PtgbSv+//aFia7IT+m0PGCRn2QPwMq0cJaCcRjDxCzxgkh0NfOl
1oHJW1+WjZEdNcsaWH+03j6wR1ALzbA0+xjEkI9MhwM3hMQ5rjhgY5l9w4xUsvWmxdr9e6oQeRNS
H7LlC2wLVf4C0ckdJt749/xP1TPTSc6ky4QrgQv+WS41t683lzWJ6M0dWdwp84X0IWvOU2veijE1
QnGzIWxcpjw1LoSdPa2QauaKBnqoSk2KypOqnYLUxAieNc0YqsTUlyrdccoJAWeda/XpOvbL/FWD
KuBzA3RKlxKWRg9y6TpFtOpGEaD69UIIjiBhWw/5L/UJctq82wt7sDlQCUXAXwNcRvQcGZzaDUkM
T/jOSYa944GA46SVlqmrN2eWTbGJW0apPuhTHLCXD5cdUzCfMiPgUGlPqCys8D74Re7hPUW7VHJJ
Z1S/NRgR2LUe3t0A8xuShhBYS+oBs1gOVgWUOu9787+Y3OwgA03J1mbLhus+/UTNNrD426HmPOKa
J+F/vlEvRrPgbWS0EfILrGFaWYKhDkBpn6cxgho3e3WAXNRx289pJZJw1+RrFNVc2Z7UdYbdoJSB
C/fMf918Kz/hPTgUZdvFc1xMfe2aL9dTJGaaStAzfcG3q17VQ14xBDnk1CjAUkpfO+n/DlG/w7yp
hz/FLUOOsa43yEE1YMyAkiiHmnFBrea25Excpuhyz64KkZ2wjLHHPh/2XCqM2mdi2IR2b3Pf1G+I
y6IifNMHD66TBdJtphzbJLHPs0rreGAUOm7wRBpqIDI6Kcyf86/GHl8m9/SNv+1v1vYgx+O9HEEF
O9iwMIV1+A7yjoFcqfP9itmIeDW/L3vwxL/pD/aeKE9Cp6pfeOu1ehjQ5FnjSWw7GeB+hkC4X8wU
9XoXKjZxtVlDr6+6FoM57LGVCZVE8Ce2aTgC2d0Q6CoxXNM8/InrYimReH7AG5XhHnCPPTsMcZog
6WoDvWol/LVn3rOkkPCKzCS8Lpg0+o+rLyyMB7mckemDMhJ9zcZMhz2x5e8+By83TAzUmHleIwCt
vNLuB2G7kcDSmqIz4p7DdAcPEYyInayEe5f3Sd7s/ycXyqp/O8yvJY+qjqiaV16XjmxtpZekQkpF
5/EvmwSEj+cUwcfv0ABgWVKuRixwG//cA9zuEOMAttR1q2C0wipzAM1VJv9JUSEN0ShlYlyrkRYG
hGgEnSZZiirm0sUQZo/Wv+HmgNa1eiLkkLm+xSFrMqv4tjBg6vkgvFYUOl670Me3+j7fU53JWT3c
XPX8zaXWNB5xxZfS5N8HehF54JFFB+9+WrGIAN8MO3Hyzz+B4LEl48/BMmpGlNMBfmwfqmIepcIJ
BDkw16xSYLGbwEHFN9NTEo8OPkVBRc8Wim7Rv8CNSUVFlKDChA3f6RtWeh8N0OktT6tl1L/6elVj
hQ74WYlw4skEXZScKkYJaoi/CpcSAJGtr31cc7f0MgShuLUk8EQxaAoEdFJmqPnyaSGs3QPw3bNi
jvYF672VnIW0qKNhLhYWBLkZ8/GlcctdnZgZSGR5MSXHUX+N7bWvHMhOiH5ki99IoKYlNNF+vQyo
SoM+BRNbIjoMrNFHt4cmDBdX39CH2Do+g0kzoNsLpZO9nQN9gPK3rIgcmd1FfrINdGuQZOB3/aIt
hCRUZBbIupfPwmZZMdyMn61P8j9jfzMftnYX09acRR9GO/q3Ldt6DrI8CXWuupmo58M7wWfJ/w45
BT1BbMXpasbB/Qp0iON2LsP2i5nRpVvnPc+bHHXUJeTbSFyrTlq+J538yk5cSdIm+q2++S17jcs1
+p5gEFkc3KhF2nEVDZ+FcuOjq92kE1QDFDY9C5jGtJqkBZloVOU9TBm2dwj5Nzs2PC7UNZP4Sufi
orkPNBQ5ivR9bRf0ws1jcfoY3oiizKRBc+NCtRa5uoQSrnBgPhjhuNWtQg2C9mtV88D6c2wH/l/D
9Rs3jan2BcJs66n57XU85ZP7OUuAXk+C6SBwx5IkIAZKFQpdKbSXZ6cESmZnVJgjUc5XzdusfvI0
HnQ6J6uxaEVQlcKg38+12/2vJMxB9+i0/CJ7RbU+xQIQ3HHclpeS+1idvEZYHXQ6QjLHSNmZ1Qw7
6oJDAztpeM99QiS8pdsI4enfsFT1mUKDA0Gx1a6ycOyctRRP/3oa8BaoaccUwGfL+9RT5Bjrz2mV
IyQg+YDTCjUk4IggavvD2nU5QZaO3jr4bPzBI0fD4x5RoI422v4JgEGciQtZBX0MPSFPxFRNW5Hc
3ZTGHZQsOX2aVeJy//1kmV8YjJIGuIRTzKC5zfO00SrlBvNLuI7J792Ifazr9rHx2yYApZBvuSEL
wt8oAtHM9Q1qT+FI30SlieKMmYMakiySZRL5kki4OKYRBnNW7e99UVhnNVbf5pO7ezFMUwwKldSj
Ks+d/lcN2L6FemAlTRMWxB1/abgfWWqr5LwmorBjBU07MDz6Qc7dLemMHlbyJJ9DjUkKjJ337f7m
+M+pp1ChaRhV9ZKv+fKOORvBSd+cqy2HdomlPTrJuGMt/W/CMQIbXn5gTFv9c+8Z1YANFeiKqM2W
I/wTkfVDsoNdxNj5ryHMMVosruEngRQQDQ+0sAcPvzML+wGoYgp5O6D3l+oWT7Rvpr7GfKN837Gy
+OdlaX71+ybDrf9u3jmA+N1FLAjMI9IdCyeA/xKSTpG3AnOzmi4hWaRhAsAGzdyjS2zvFY+F9sVa
d8UV/hFP/gK8hVKeu+Yh5XZemCnJgM0bHhURzSDXXducCM7J4ZXW6/YKtB2gRRlMPU9njFmXP80A
pfBo6b/gtAJ1B2tzK9hFs2DoKBKPnWKWI3LI6xL2FgHWaEdGtsEQHQfCP9gzOXPdoHQHqDwJBMVM
DFvjZt22MfOhJKENyhiNSRaF5G+po+0mIMYSKWAQCRFgFotCxwyRNYvOoHQuQNlBPhG4w6txR1E1
R/gG3jxRcU1Dr6gqGjeuuJEYbAMe7Q9D+Jo6utDF3i8B4T8r2ptm49unTB3E3NDLXrrcJK6vZoo8
TSXPUZnQZGnJOekHoXjVA5r54nzZJMPNhzBrfm/jBIm/wwBZSOVcfKhP1R1Fa3U5eCkhSWMVqvS+
XSfP057bT1Ytk2l73+hFBcggjYXX2ynhoos4fPBin14GxKaFbkCvuKMH/nhtdyElQg5/UmI7S4LM
nckCYMQgrhrOI112UxVi3l3QpXoTSKbHm2s4vBhzmrQVx/3C3L9ueyyv9W/WZFgHFPxwrqHKV/kD
1wHcBCjI9lO4/u5s+DGUvR0bcQFPVIzHkY/TXMXjriiIvkhKGWCO5OOTWgfKSykhHm7hXuWb4e3R
3vtbHy53VmzO2VHyzNk0MlfB9oyChLxyrJKF6sIGu+OuFOCoUMbrhaDxarzcPpCNTJm1iaWvmGmG
iUH+hQSpS4vHlCBsAxS5PKXhcH/ZFqa78GQJo2jiFYsEhX+NTev3JEH+b7COJuaFyjHKUnOwnjFj
RdGmfJSoVZdy4T6qrTTFQs9n5LJPYF+TBtp7dFyJ9MqEVklR7o4kIZrVkEnXlrInX3JCA+ris5Ss
XGDN4CgkT83wri8qdpZ1QUBmhQXu+nPe+eRHpLQQEpTNtDseHRgWZIfFeiNZRe8LsjxrpX5L9eJi
Kjg1F+Z+r3iD81kiiQSjP9MODLbNLzBZ1Mf1XBqR2qabrA6gLufo2EjzyuXaP0t4gnVi1uxc3ugS
yj8e1fRdqLMygo+lCtG1kcQF7Kxc4g82mk1hcltKbn3oF5ogEinlpKKBThbQyiQDtgMdOqO/2aPm
nouHqBs9kAyQGxvMPOV8/PF0rtNu+wxKZCLLVhl5VmsxQ/IcRCxJrLjZWSZv6zKFhXUsldz6ZUtd
lmkFzSY3T9V/hJcQIzTB2ZZhveTEhnrHaXveujy2/oCoe/NIr56Dz9UVipKMeKzUCJ6CLYT4Fkvi
eR07HL3yNbJXanTgwzObgg3xCZ3hBZvqbFZqwx38F7miF1GQSVNP1B7smTpgC04T+7S5gIxnfxVb
JlC7NV9g/bHnkcOi6ykSAAHVXORYmnMj9132GBkuvgpS0KaJZ+qNXrtkncOXQmUBwH2c1Ir9Ohyd
Fud3Lnca5G3fMEa300RM9JnPUuFjT90DH9McUzI+VyT8QGyveA37lzLXMs66ggrdUzScYaYusMpJ
R/56qCSJqtZG7ZK+tUCPyvbABarvp2OTNBA2jT8OTmfA7I00WiwTn8oh/EDQCcPzvLAgRaUMO1VK
/lAJKMSRNRgxoMPgBxr1qlIq841bgvDb0reVB8l0sivNDJCsWi+AXvHRNDyUuot9At0nqNN2YpR/
oC0W6hZFYKbxv+MBeWlAc2QxXxj5Mb1gpJHLe+WvSYfIW8CSUEmTWmQlIirJzgyWGsKD7qil6gIj
Y8bWT3YKqK6xBg0VtU7JEsudA0Llr6RTyee7VmeGcLUzLS9H3Pyt903gnZNiWNz5jZGfcoYDwtjo
eDQZAyNtY01CM3FYN0X0/humCfN4U8g7DZMHN9zuIyCPWUUj7pcOJAQVwMHzERr6dz38SwvGULAt
XsWBlYA51+JvuFA240c5qMwALVN2ySqoq6p7CqwF0ki04oHgDmau0AorhBKIxKLxEPnO5xshEg0V
vDcpCOi1ne3BSMoo6813scJLRGByH0PnRd3RDU+yvojEVS0KzQ82BwXrXLsCVT51VEqURfBC8o/o
yTgxGsIvEqHpXRv9w6exlMef7UoaPCAydjI/cv8YUxtOJK3lGkxMFoYF2S4mywxbZFE2lJ80b3IG
o0a6QjxfMj04lGxSUwW78YLKkSnLgRV05A3UpUOuT3eCIa4f4x1NA8TMvVgMg1OMMiybYilkAZOl
iwHN6hr72oH0fRN4qnHgaMJkULZNOAQ1gXCFYoQUwNmxkV8g0PyYzcrZ2vqKpO0aBgOHW+r1ZB+M
uFaMv/UIGDCDd3RxbEUdA3p9SFppwg/D2Bv1OmUTPQLdc6AK9lxPWMqK8M0vn5TibBvOGyOhs5vI
K4q9D5KKr+yQ6GcvKb68P0vx2GWl1CDQLrUBiTp1dgSff5Jjj/NyRP5sAfF/QWkOn6kpXsYJ5ALe
JmfuYVjg/ZdcIp5dJmlqdQ1pyd/V2A9oOjcjfdlILKd/w0tDdtSV/iCpk8U5D3zS2X0AzvQXszJV
sQSSqYvjt86M7j1F5b+jVBgQ+DkJ19ecBL6J77psCBMOsuaZ7soGjXMGvx3DpuOZwF4es+FXP7sr
cYhlm3P2xuD5reT4vtzPn6OoSVsRdVJdGPH4TdI4cx3U93Q/NrI2jGfjwhed5kH4OBz+bs6sNK77
4zPMh08CDNVWWJCwQbSh+XtaqcTNUO2xsjAPfU/Z5CFAVXbRrsFbKSE17NKH/H78z83em0k0yeEa
9ab/a2LxNchC6PpuIgAoXm/OBOxQIqnPIv72JxbNfH9iYU92IGqYI8a8xcENlpLXt3D71FCjnfwB
s88fQX9tmDyMLsd/8BzwId3FVussOd2jqRtJWmZ9SxAOMh2ZHWp9oKg9ZO/2oVnOlZRYeh7hzcuE
ZiujKkMECNqGm2nyJTdp68e9Cusn98lArDdD/HufXEptyM9Ls4x2wG6CCkEHIPMqmBx2Z29kyT6h
SpMZKBGVyGnn1BImnqbjj/JiNddoo2lrKP2aMfXdJ/SqVQnrrmaWSqoNrGv9n5bmxJE//7GZ9Ru1
5SH/t3T2DmW2nAmtP/spcwW8NpxQ84/0MYezVtp8rRUeTLA8joFnWAd3EZSIqOP9OSk4v3eOTGeD
wseHzj1RtQhea2o/TaKteuvQR79jTXUhEEb9+9QC/Gi2vTFZGNXT72zKaxCbLyWdCAaPHON2ScOS
pglF+57Jmns31Boj0Ui0mwU5awP0W9br9o+n40ruOK6SvosSzMPUMDwg+MLWD0sAEdNBkRU1PNpf
AUf8U0M7PrgteGlQ5F3oe7pZjrBoZK9hYWlKIZOwC5CEMBiQs6CjXai2Xgyh5Af2RwrPN0jXMCVJ
9x7oJT1dz0d7cS+CXiozWd/wW0fd1lD9Is6DOI5Jz1iNdtvmR6EZNd4pVRAsR4SfgiYGkRC/r/DX
sFZw4njkxMRmZklZ33BVzEzaRsnxqDH/HqgW6PWR3TY83Q9KLPKCYLSbbNdarjDOYtHz1qCs5qn5
5sGUQQ0tOtckKiEaA1pMUJ0Yr2XYnU+3E1BtkrWUqlhBOJ+HdMYeqvT+aWYsLkWl1UxNAqgjPd8b
h1lAFQa+PtPK2LUg8vcjEyFaBV9LYSUsFv+bTZLjnAOYZ/EDbA1ZZKxikD0s1+7CLE0V4Xx7xaAw
035PiGjlGT59Gq0BEcSkbQ0fFu58x4/DVPn/abl+fPMzGsuudKUNP4/YBi9rEz4MxnFhJjD1NWxW
HqxLRDwY1DVTAX/4sTjgr+hXiWP4XZmuLP91lxQ7JM45ss3hU2vQ/A2HVv32SKQlLRJgZF4Nw+Rv
Gf4Anf4ZRt3SstKX4Hzegik5PVzRT4f+CqjS2kLddIyBBYuEbKtfNdwGnQxO3/8iazYThaRo+7LB
SEoojEMzVYPNUoJxpp1GyWSmR9Gytc7oPx+7JqQyFrBEvX0OU5KlKjjE4EPv0jLBxkqiAKY/OSO5
mCEYTp/g66jlCpKNDXA3otVUPh7jnwWKcyLz7uP7F4lWJIdN54Z9ics2SNDHI/NdHhC3Mn6+emXI
WSanQwCPW4wX6BdpvCObIVuWQw/wUBXnaTUdmEBf3wMD4OkdZTac/mRJkl8j4peRoFZuFs47XvBm
UOqyIs9cAEPCUsWLzO3dsaiyCRus118A7/QX0nwx8hzRuRBntTQfr20efd0FIuXGZm6te8cM0jjn
h/xWCGczku1mb5ByErY1SNDh66hqWFfF/qh+CJxzPZpRg7AmrSGznh3AVNP13ENjTQ/OC+xFeHLd
vh6ePZRhPHh+SBDhL/bfIpLvO0lEzMlioD9r7SDZ2J78sd1y4qKPVM/U0XFLjzFX5P5mA2ZhBz8h
WuSRWjUnOqyR1Z0El6MErJGG0yUF+3NqnSVrsOoFTNiZs4V4haazHA9awobneBwjAsmtVDknDbur
MhVXcLUwtv8Khifsrfl4unJ1zEke55vBbbVlGuDmNMzl3YHxSht3ecJ3eSngydkCDN1buYWLAgqm
oRe18Y01xek7igzZrmP6J9twMWaEPDCW+j2qa0eLJZ8+3Tdun3GhX/jIDElWfhNytq7eI1YYclhP
WvK8ZFFLNUlZlJHEQdL6cVMmSqjTkDkeGwnhKvHh5n6JybaxLpcoxhDTgwygAb3+OwKeLToU+A/h
PscfM0vc9HUhlqQfd2QRYTf7gndkdMkgc5LEaTb9/flux+AEv3mepTh0Q+0sHKVM0jGl1bk3cFr+
963bvuErwxTZqZP0Pyfw+ubi04ALmOVPQncQM60ZIMfu3911TDhxB3xaQkNYwVNLUdIVy3076DhT
HkfX8Df2Q4l7f1WtpyrB3UKxd17kA6vbgjLX4hZHPyxW6PQ7gfzeVf2zsMEno8kpzdmQd8+C6NKO
Lo4FEpak+T2x9UOABha5zqJpqHc03kflPB2c1XVwS3kJ57Hg1tYHJRPD2gUPMDvVse9dyvJVgfYP
KMHGvRrYx+cL1ygzj2tJc3K1Pq+yLctimqSOR7maFzTkHZEoUfpEtF2LcBeqYZKHfS5+LUHEGssR
GMUmL9YUmltGReUGUcmkhqL/JP4isGWqUsThXw0qqK32TwXVDhWu0euaKPRm3QUiRE/OWidopqYs
OnVPt9n0RvpaTf2M0c5QW2JneLv+TuzSdM6WQg1YmPYQg+BBZUkzEQ7VSlGSGLU5rJ1lwdnLejPQ
/ZDZe4A3l+UJuJ/5/s+EK0PIR6zM8QsK1GveyfG8lNFl7vJdWozRROO7/qBv0eKxRcUkdmYQhqUN
v+JEbqxeCemZNhWI6LD29KHsJ5SKLQcaPXgbRIGGwOe937IyJWNJOP6Zmx9P3VWOysoiYdQ4GfyT
JrwfhULJEzYfI+0+nfQz/QidmTy6XHVpr2UeX5j6QWY+8rKPmJ4QrKIixNKdHZ/cdA77OhQsrT6k
c5jddgzqOmnKyKn2y5kdMdG2LnLUTpJf5LQzhOL2Dlmb1OHYv/TBPCpb3vi9k+KbXY9YLF4azy3m
PJ/w22zjtoDAeWJPh/RZ5u+coa1ftIpeZud1qVoQBSVNPe1ZPicNihg5Zv6QYnVFrtgKxlh9y4Jk
HakuyPCv8juEN4ZapeFRNG97w+z8LDlQ+4WwTUqB/oiiZrlx0SkB3JxS5YIGwmKjMJSoB1rBTE96
DA+InJWAguzhBrMctAO9fiyE2Ake+960GZ0TxlXOreG2kHgRyhLthbiSigDTAuTfkjZZkvZY97QK
e3dxXtFC4Ah9OFkYjsgGmzjD37E6LDVLAuM75eSiCNsuooIWjBeEobFdmX61JIvcltKpQAmNcSDI
P3EXPKTAbVlnnSKlUHZbW7gNzkTwsWt3j4vmZikBEosDisckM1nBFa1adVPDdQ50R015VsNKAvlg
TTNzvKeBWuRgiPUw4uV9IqVEGxAVrYOfGuMNPqyWtQrBdG8rlAPOFUNGufqfcsJYr9ELJNWB4Yc8
Ihe7FxrzlBWqiGhqcu4L+kzpkOp6TH72pv4sQ0T5KE63P82MzRUzN245dCUF3/HL0wdXn7ZXPEby
MkkyPWU9ld7oBrmo0yfgZ3EQlSeeRF9O3ubrVtRaa8EcJpCOJLPIp3L7ocX9dZNYs8gDOuFt4lrd
TxF30xGjnJhINVUb1kmzscGs0LfltvPghDX9GkdcJYnbcVfmgmBh3BryFQt7xnHTEN/bPWm9eebi
UpPVCG3yi1IWgVDlFhlJdcJFoU4hj4/UDvNosu4KR+fmbpSfjtu7uAvlb9neU28uUn69f84WZlNy
ODZMEQsb6X4CgLtBee3bXAoEC9xI43e0GaVj7cpwcQNyUx72FyOfh0EGgkagvXyCzixeCFavljKG
lB4oqYZsppQ05nrf8q1xWBJk6PjC7ozvNzF6BjDVnRiN9L3zP81Vb2ngBlNIQBFjF5x81oaY0R+F
EoplfrN8nnnNb2bw2HsuimWWEd7YwZiomYlb29l5e49iYr6CGCFJeqVYKx19nAg7uhW3id2BrYxC
Av932DgNO3AeaFN/1gQ8+x5pSXrXQG2a87qZZmwxaNSS9yDFhNwvLSVFkTUjSCJDk5CEhkay+Vme
KzLm4+7ViyAHGwdIIaxQa9a8mrdpuzWM9LRgohpaUkTS774uTs1xYFL3yRTY0NwTBdBLZA85PN0g
MNGZUlcVGbVru6uz1VphMI9iieJG3FCZpzx2yXppG0t2YBY/x+q1GLHtcPZub5n6G35ZHFPQfws5
p+BiyFX/P4YRw/2YnT2nopb7xAamUEyBp0unyGwFJIN7eaUB6ngyFoVQiqVNN/wyhAF0ZLC90xZQ
nX6YmCi4wlUIbtXXIzOrzs5ayq/0cdDHe22S+ulbqpRBGyo2b1uOQcGPd6iYXM7GlhYbco6D4mvz
BjuyoKb7iOutaTJwuBxuRe9jbi5ycgDzJQc6XDXqrIlupzx1VdXmt7jdEhDHdE+iqhKo7l+1HpEJ
5mHpTv5jS/CdkDE+syOR1xzAgKTzQgugeSSDL9BtOwwdRlTBxmzFOmAS5gll844Ww46J+wjBzZVu
RQ25ILEXVHpbxfpVcbFE2MZOVE1/e0+OyhAuOztBelXx9W+nxjTmlOJq5Co/e5G4DFQV/n5Nsonp
wRc7/6/1wnu9f/Vo4730Py4fXHidor0/BTG/Hl659NGBH2ynfM2ECmpoaxFqcVIOP0N9vnN04sAG
gaELgSTCqjzY6Qwna94dkKpjdDoA03/iYcjKbEVi6daawf+c3NsHPkDCDKDCxP6n/6061CHr8ahL
/9gsfnrEa0X000voqo5PpR8hysEcq66v9ujwdhopozyz55Tud9IRQxBkXOKAJvHN8utOr85HJ5dR
qElmYKlwyKmNQoMWe2q+1oXF3njv/I0x485XKSijM7oIdhriAEV5STwphvU0V7EaZSDBuO83UU+N
xzALABwef5DXLAka4UnkirjcBCP3tZwXnoYphDQcmF5HoLUpaUgLEk+pNLJdbzcunR5frxkSpJcd
rD0TMH3n9cE6eL/HAYxgNjEZCWdCP8SvYTFSVlss/oaoaI8KVLoMqtSPZokMZ04ykLg3zhqDqdFg
1uZY03jeDOdeJzYUWSwCpNISHDzms0Xs8jkGU9XXnpx1zkrpQBI8iPRStE5/9bS8Mx5+Zjkyy+KC
g3W9rCV9tvYbyGke+uiEhBvDtqoGg09MMULxckyG9ER655FCeek73ZDLpfDU0dx6Be6Km+t3rQr/
hG9C4foQZwE0axCZs0i73prW3jrqCuFJ8uWNHT04lBdjgMao5wNTb/AaVCgdVKRPHAW1+46C0YmV
jIDA5XNXcKWGYRmACgBeGLnssxm+a5zIwNyIAaYcnMU3RLZeiGTs7UoK+Rg0dp/dtIC6OESTDvQn
sjGlsga3qa0zlGK47jmKSxxgPv+3lQb1Md8Rh4qxLLS2SFKNZ6VWAtJwo6NlBVWrKHavPEO4tOd6
J+nK3Vr75COqcXrJUd6xEDoAq1lTgE/zZipzEGES9EfUl/Vor6A95Cj5sep1pV+zp2SRyzx2qqU/
7W+8UWuJFPxhAK2/PbcUYPFhRt0gnPEXn1br7JYadYVNo4Ku7AtV/z7v9nO8rg+MFRkbNeyGbPnc
6UIVrXONR1ujFCUn5KFn4tW1H1C/PVJq2cEqJH/APRX/LWG3tmvUwWKp8hiBO64G/KY4bdRdYxcQ
HVvd7ht97cJcR8dRohXZcdTPoaOMQB7Ipj51mlUmUkIwfDEnJA/gS8zS8XL9Wn2Ea0iBaCuRcPzx
r0rKA9AvmPlSr1npC41358u+ubRkSv71aRufYDmJfwCGO7SwdPY3Y2yA+D0UVf8ZYJm6qvCe6oE3
ypQOhBMsIrKJFZU+clRg6N72/qbUkBg10UQlU65FrqJP8lFttuLRqEXSwxc+ucfTjQLvngYT3qe1
X7kt5GhF0Anm8K6BFTWRwvlX/4+5wBzqTUOzPBWCCIQUfmyN1VhOSqZ5U2uLf3iDsIrN+malMHPg
CO1ouQhIGsJXU5yFs+djtB8Xokixl7Z09z1IHCHick7xhq6pXirHnEc2jjOJZT1oAUcSRSI4fbw0
n4eIPKB9R7fKOZkBoB85H56gDFPSwFfeg/ag8zhzwlwHfI+eZgTLMDxRIsSF6amgT1mszvmWw93k
rzTO2VJI+MNYtqZLl/LMpYUMDf6y542sIb/7UoZwBlUzLm3fapoDxz3BGSzYCCsf+1UAWiiMH3yl
ttcXXhD7P7S0teFxjyBl2sjnV1MbBplobSGNt/CxdLA5P3FgVGluWo0MKgbrki9UmcPKWd+kAoYm
0AZ6JJujXrSMp1ibN3vCPO02W7fVV1sKaiOvD8aAvlx5YVHtP4OObtyEvf6YyumHsFMS3+H6VSLk
NoJsBsVC1mOLckVtg+o0swMWobTcCfUJYe3gN0HQMknn1m1+Z35pEu6ImqWjuM+JkWMWYNdb8qOW
Dzkovpqx551m1oGU3mmDGIVWAwSxHPJwvnFyrOI5G00kYhIHArGjN3JJHtRa48YF+Sm9zniFRnVv
GlhOv+p0HD7/INFkosErktdd4RatCrdGQIamlFphVTiVvoh2bJ8zJ8TniBY+ipE4ITnc7y5bUnN6
jZ4PQjbMbqJOXeGOB8c2BzrliVEATSIJwxhsuCHPXmX7kui+EZ4yK70aZMyI050JVl9rqBmXOWl/
J7IjYwaa73XvT5jPpzsBMNs9J7DtF2c9o/nFfAdmpug3/r0yy7Oi+IsVFfdHufxUXXOV2gV9lxAV
aE7sVhXztuV4P5VhrFhV4qbP9hUEg2zGNAlWGcKdZcv3RMEdN+EAAziYhg1NdrpApmCt80iR5+y3
QvwBfRBDR00YUVRWE03OSqvlGxWpFO06fd3tRVCqjiTKrg1Lx0RZShfhQf/EKPb/V1DWaFmT9scy
DyDcwO2l6D2sxzcqs09viWIr4AOwIo1kOTXY0vfS/kVCdWOAr/EekEmFWo1Telaa3CEjKKi8UTOc
EHPkFaPj7QgHhriO1X1gNpu/8ZJRdpwIQ43nyZm4Q5T3DouXzz0HhXFZ5EOuBzU7QUsUlsX8B103
cyA/MRRHoj7tHZ92sgeBA19k0WzdVlxiIWHXbkWkWw8VPe6wpdr9CZ0J8aFZFTRwaGYtCVWHHGIV
5I0NEaGXv+P8sNJl5LcEQJmyRq+dJY48C5XHd2KrrFsKklkTnrIn7kfgSopBo8p/vGpfMWkGxWCt
X4rgUzs8fCTeZpDd0i8a7H0f0yXtBO1TXisyqYIFiPPlVD7zi0l/O2GDziVW8c4PyOkX8qFJDQoG
NneJPKWszPliZCN64wY8mEU7JgwlJel0FpZreiutiNYZnl1r5q/8c48tygBG+OBPw+4BIOXK0xL9
MSbG1DjyZord1w7NBeRhLZl74r++tPr9cQrcAABjjWhVmfa3DbU9HE0P7ELWMRtnpfMbEcdOsGSd
Eg2M+7+i4cfONrva/YEZCuzVadIII/fFBz00tjOX3hH6DDVViWQX/H6qF7uE81rOkPLkaa0im2es
THHLgcYJGRdYXB/NzwkblcMeC5WbA32K3XC8gAISv1zVgacO7tjVFf5eTyPDA11580rXn36amNbs
vKYaTSCqLaEPnl5z8tqVm9GcLsgVEC7gzR70l99kxLHTnKsWU+58JefP8I4AlYRouZvT5X3Mv0B7
dDHLFdZ3bOZEVjZ/iy7RIk+yo3dOU0EeHpN/OQT8/17XXOTSAj+MpeJUkLbs+ERspb1disJT3Eqm
LE0FJWaxJNbGUm5+OK2IESrbxDV0PpbCo6V6xWdCMbVlNQ9eQylT4zbwahpMPjIxHZDpGKdS8F0h
q6VKnIlHKG16TQsVegmzhTqKQx73vU58x96Q9oC9T2MXMxFnMPZg3HAEOOAeV8OQa9jGxyGoNNgP
bheKEQ1sDcETW3cbvzbCrTlNiV1pzlFMb07Svx3X6Z4gxyfsa2yOiFDHWEu7kIB2gk9sgBEKNYEB
jUfalJDe1QYXGJNHzlCoVHqjZNEijbk4AUps5GaAaD0TyXhpsY6rWknq7ZR5Hz2RVjm7UeddH+jY
PJEu1HoIKXxRHiSDuMpW8zhjOAaDmPzRwSLTQTcnCzUepI4SlYrq6Q6F7snlu9HCzE1Mw8LulF3o
q9MYKWfErPyXy7bocMSG6liFn1ju7MVZiMv8CqbV72s24GImE1wm8PrluoxuYCVEy61xl7tavKwE
jTnaVKfco3eLbb/5fF30+sqKo4k1RLuWa86tPIHmYWbcQorGPFLNKmgIGcq3aAotSec7PoQVZ49J
xusVmpQMqoUhk+eOk8vHUsIH+rtW9IKQF1E3VH4rWfiLziQp1ALbCa/RZVrvcWz802jbVkGK5qaT
ClbTQg5Yi/+v8FKUGimnUbUOXIdIgd4vcmvZw7WGKnOvJOf7L71ITu4YBN7NIHAVmZkVbVPpZj9b
uZEg5WCf+N147SJ0k4Uy1zbhCU1SgiSrtu7nM9IP6wBglv+vWKFSiuvICuLWIDm86S7Qd2I8rFnI
vKATSDRhs7OQ7KC2ZejkY5Dui3OvK+nSrP+GAdS+OEwGb0f31UfVZDxb8hkGfiBBKuZbxDJHPlT2
iI3ymzh5mP3arIzv61iaN9BdaMGlPHg/++Q/GbAFSVdkWVcj0b5JKlQoQaoxEdXCzSWcDqLbDOO2
ClhecaGcBDwrHWGCw0ABlLPmj0K8zribubnkxUejclCz1qdrEIaXKWjW2Keyjd61wt3xfrJT8qeQ
MSNXuGur2UnBv107RfpAPwJnu8jaYbMpv+aAYTa3K+wOcWeDLTYxCqBM0rKEQYuJk4D11LrMk0sL
y3aCsKaWgVnWBnqRmZc69LYYcpS5lWlu9greYMyShE1Pfvq0wtgCwT4bF1O2oDVHo1Silp5CGt8L
Tkf/OeuwDIpz4hOaMg8t+cmz2J5ABW7pyNPKchT73UF3LNWabSn+i2unOd+YR7zYpvInw+HnRq9q
QoXUMhlJmaR0R74HQYOabpSj5i+lLX1bV/fqPxqxJulLbskdFbWa9k41Jg6YO01fH31pAvVv2JmR
HohZvi3iBcwktRxji47ugffmMighRWkEF+9fSdesvQpM9InTB2joUBgjP5+I6ypffDdQGHsS/oCB
YtUM3Syo4DsSXlD3fKOnGrju3i9MC/2bP+NlJnxyQWrPy0Pgh7RQJzNYfjcV55MERf/OO1BZ9TiC
lO6sfPlXDJZlHLPF6DU68Wfyt7iaLmhN1uI3feH6eX/mvv/CgI7Ul35eAo8IhnYvKMIgPA6M/Aic
TrGrinyptmX3vDARbm77+/q8k1hF8jVOeZRhLmjp2CRUudxz4wn10reFMV94sFKGgIz/GA+6JM7B
O0VE5jKI0azD0OJ1HPQeNxpq7dGsveUAv26uAWJB3qSgUc+niAfexUtSt08nMFYC3z0AH++RRw7U
Ty5frmXWKqqbH90BZAONYEGJBB/vgA5nfSZq+iUTNGLxNztNUdh1ERiwjqqAcgEm2rvcktuUGVYb
v4lWY+7spcFTnNIxrAjqfJW3ApicVjn6OfP6EAbcsLODYMp/nYOiTVSsMhLT6wvp1/uPGJoP5wzm
RKFiUfhYh+gKwSXSVtK0FLkfyv6nlyrwskgPcTw+G/wlJJhyw/i5vkQFxmP/TN75TkgLxBXUDIn+
IeSUahxAxepYSdd9m4fqzhpNMqE+VyM9fG8Zg9cXX4V6P3B1k4Nzemn6zuIdfQLgPro6oCQ928lP
/a0yta2pV3FPNlvrtzunYhg+ZVV4yUbAE3nx4P6h1lEr/skDGwaoAhsmyqdyy9Qs1gX+EWiIG7yk
akC487jwrBT5fYN1Bfizgz+K8Oudn1m7JmxVaLnHLUH2YndmybXHKnnYHRRlSdME6D2xAofk8lBv
rmai+hcYLa2vfiN0AWdCm6xNMQfIWyGuENJNGuHjKIISIn8PSdFBHWDuMelvoufbg8DZ+HoW5Nik
8z6vQkAQfBVSNZHtQ1uBVwoxIhzIG8WiNlHoj8TnZ+hmcGwT/B8iB2a/qnAPmBRzH8knEsQfGzGp
QqYeG50OTNsrOhjkgv/hJDfb/f00pHyayVrBRywvxTM3C5TAfYAe41V9w+vGn5XVfD1SHPGqeQ7t
O62Egmn5gKwTz2P1W3XXAG525CjPE0peYo+fZZhRCs3bMMMaWhDIh+tDOB7iKOpaE9QmT88iaIGp
GhoJ2bzSbftq/AnT6wpJ7bLecLHxyygp9LWRpJKEA+4KdRvDaI88T+XjQUbySamVz04norgV/k4z
cHAIP6V7JRxQ2hU2IM5ydpftZtKDRRlQxwIvE48oXdBxXXZnyx1EUVK/1LQEB3rmk3Vrs+N6QkeS
SoXPPvPjc66f1eFJdUqkvS+lMgNMdOdjfi/LemJFqqcMC/PMZdKUykubRw4tiY1d0s9IedjRuxY3
DP00StEJXaZ7mSoeNsK/LspTlpclnmks0ApaVn/py67qJG0nWkXmL+vJ8iMxggWnu2Rl6SXL1EYH
fYOgZE2MJFD3B9HRIeJ/KYot9ik/t935/OdVdcmFNLulaHZca40epW2UH8r9uZfuzADLVCjIUz/r
P1C/Uu9AnWJ+4NqeHwYDWQ36+TZaJ2OZYg0r7+Qp5TGyaBIqYkX3TGrjqd2WxlDV1AkT34WtoIPR
dktmao2nL66RQAwsYiScKml+gv6/DvUW5xwfFmbE01IWys0/EmrvU5TP85c520Amv4R4WaNE3uni
P6YBouYJmGiD+V2uKrOgwMa0CvfMEP6z7ZZHP7gNWKgSc2f6+EP8nlOIdcXjl1S/lMqcB/M1uQtA
FyYpo57EPvsskwZFQTgl3iTaypxWrsUj+r+o4digPrrueo2A/Am5TqMqPQ8AKTm+pBy1Q7kw+zEZ
stRRq7NnS4olMmmFXVUcNrDYTYRuAsy09f5pR3Or7RDL/e90pzTij9FVoKWtU2BLrr9g3irdq/Sg
x/EWEIJvlweMwHounOtE6Apaji3LS7eKGQfzuxo6HbJVFC6uR0fqTyxDkYvqX6fvrPsBRHnYHb9P
8llFcMUJCki5CS9SM7NPF/ikXD9MVJt9Qqxuum7GH8tgbd1H5AAPXBmVrdUYOWR7trDfhqpOZqj4
PlPiHW7liNpeR8BfoTPX4pJmCsWuedqkSRedWSuIpITPrnhkldee6Ae5g7Etg21MAWYgw6audn9w
sv4cLTKPAyCGJJ9vdSPFICZlMVwPBmanlmqVhcZNDtAEmazAVEzEDnZlyM7oBrFYSwZdJJ7+/pIh
E2NsbYJsPynb9TErcRrSUAychZW9Re/nmdGic9yQY9wj1xqK1SkSXbU3XDj4NUgxvtD5koZC1XUx
z4Y5EOeTBAe9z094asU4nJoskcIRN+SC3xRisPbfBHbA2upYhqTW62Qtozb30TVtU+fL+oEIx+fw
XpUg+FrcbuNOwEXnwK49C3zaeshRpn5KG9eyX8+M6bhFFiu65luQWBbxJnGsPhlHYOd4gPwbkjaX
7QcnaZvBClrA0VCoVQiwoW8omRuja3bZ3mSGiFs4eMwxLfNxEgMxM6+a2KpDqHQ7jHrIZz2oUkVX
hr0OGkHn01HDNwEhORS4MDM3V6Ekdx6e7R4QZUhtglSFI3OBTN5FRaAngViv/Yf56XSf+hq0WkDa
aOZlrEjyqEmMUErfF3A4lEgXb2ffceSLNpsSuDGGPNtEyzjPIjG0ftxvudN2LVEpyL2IXvmjO9rd
10bU05ssldh8xTNZEMFTxUBsOcS7WVqSDIG0kL2XTDnS6NHGMp1wBk7A7vw0hRuG97Komg6xZ/Fg
DyAFvnncH9YsX5TV2bTBCXlKVGqicOXhw6SfNyV5CikvubYwi5SDA08HhaPyVLmk48YLhwF2fNZ9
cyYzjUDC6ihDA8scHb0Y0FSnfA/yG4PL8xuJWlcyrSXK//IcPgdwYOzpkprK/kZ4e8fcT380WAXj
uF0s0/GxyFoWMrioFh8M+zP1EHK/jbdE6Ywupi8dRyHK9nYvUUMAezVG1lvBRSlnEH5C0mKuHg7I
YE+aP9hz0PL7/T8F5L7LDOIxeRdddAVDEkEFJ3e8ZCv27VUuplM044tGfAZW7X7lVjrd+7GFHtvc
P4/tAzfee9w9jAhlg4Pu6+7sisXf1MzNM4gz0dIUE0Bh2dap6WlpmrX5GXogLKKPmA4HzV7e0hKM
P0WOVrSR4oniwvRBS34dCU0x3/3vat79bkAYz1yH760pf2f5EbcuCKP9ZDIujsdnTX2HsPTSujWN
DL81Xd0bhTJwkL1iDSIQfKoAlQLmkZYSwy0+Uu8R/G17VFCTr876U3VYej7uI4cZrVYMbp6f9+tr
ZcOcZyQSnNERfdyuiRb0cuaQc2q8bOhVpuTfxULynVtcwCIQgm4V/FiFLmKHLFxQAzYiyVnJWVEb
D0TrE4Kx5vbq5PRW/iNx6AfMOIUSzRGGBPYSI0e4++3xu1uH/xnK2RJUe7H3/+bZHLPEI4BQdqN5
O5Ol7Wgn8E40dZCVht/xX7lrZC/RREVulnUJOZNCxq28bV41mEugoQJBRR1rjgag89gmng0GUYT/
pzuk6YKMfJx0h77Es1TRDkpf4R+d0iP63CXWSANODnzaNlmVYvDIAEkD+h3kCojbXMT7eUOKBHgv
ONCpMrT44GCG1tUh+FDLD/1ZXOB0E7DeqOj56sF/Oxtd1fcMbWSDVH7OT9/T+C1kYJ8rgv1gKZ2j
NRrmkwAOsZPBo8QgI76IYqdGKJuoz85cI1cFPxv84xEkU4Y2VxAMoQL3v72KXziMVx7sOW+DOVbz
5cZGLL1YUI2LW/iUn8VRF5tl4KgM4DM1JZRRyYsafyJ37oibKWZLWIlLKBpKFJiy8gkYq9QC3Xix
y45Tm6vNiTac3fu4JaLFCcBc2XGUiDL/EEMIexnV2J1lfZ5/JLBo2j+li0qVt0d12Ma4hYlZgJ3d
9W4v8M7VCfzVb5qgK+v/b80JkmU+sEg2DFi/chyaGw/NV5xXx35xUa9c712C6e0tlh1DZgmASjiW
s+Cgok/jHhlrqOB08BB3M1+t46HAsOyY1EK0Ln5+dqgBZgd9BFUYtRJwbpNseunytpp0Ye3qPu3s
aJ9fxR4HCo5Stt81gnrc2D5bKxmjMpOs5UrhqunehxF51wUXSPZDRaFoS/qCF6QUSgW8Lecc7u76
bi9OMDPIvMgqqbO4umYcOaso73jkvdU4SHT3LJLg20RjPfpl2FLL8kL4qqFaIYPPu30rMI+QBv1c
eDdHXPAa41wYjK2PpDg+3vkfZOHj1zszYlNN1QjX87QD4cgiYX1yDEta5reIHL5H772TQMvDWFZ0
U0GDNRvVN/cPSy/8CbjMS+nHjBR7F6ym4W4Luuas8sXVGZz3D9Ye6s0NEj4tCe5tww9Am8lMJ8WX
lol1KCKtEMtYfdq6zw6XLi3xZVXFHEVE5Gbq8/DVNMCM2p/scGPjookVgP2rsvLruPgk2/lVPfiw
t3iSFyl284UDXoR/2xfkfw7+PsD7RJK/QH7lORL8/jjouQmFPAIc33IWbcfsu+JHOWeNWORUaIoL
fu2pD6xYyIGLwzUEbzfCb0wLyL2kpLyYAIbPTA3pm07VwkjzLnh01XW7Up5MgVzxMxKCudh/WD63
6dUznMbReqcW8JWRm3aEQVWG5RMJZobTP87m0j7BOm5YXmSGxZ33sSWUMbEZTz5p+UFZmD4iNgiY
SoofuiI23BS6+gbqTo5K2E81lw4A2agt9QwfLVKYfTfs5r8vRlHJ/6TdyIGt5svye0kYe4sw4bQN
rcrWMmnYHFaTTmHB4h5zJjSaMwnt/WvxnQg0Jul5wCTsV1ARkVEzc1c+1EJOz9jiMYKcVdUW0y7a
sf+g4PlZZNgphauFXiUNs2L+59gaosVsfSCWN7Ccli0GWe7yZ1+u8WVykTZJLSiCcuCstpRfa2XP
gN44RlOJXdBNeg954QuNO7tG7lb5VdUBWR43NJZjgQSozlOxx/KpUGQ970DVYR45kfghr4YM8Ood
geIMZCMZk2K8hlf6qGeugJsNIBp/jtSkWrtnpDL61WF9ke9WnJBe1Zpbc5vgCAgfDll7kQuKtned
DYBwqqPw9Bk3pWtjlsR+seBApiq0Rrn7XNyZoPvfGyGMYl67/38SMMZHw42ftyTE44vlHc31+QDS
px9zdTaY/8eBUZFONLdxsTHZT2SwaggB2XwS0ahxbxPBp6r8Th8ezsbb3/BYzOJaM6zXC2TbE74b
f9d3Nh2O1yCO7Fc5lH8abEcn1BhyK8nxFLpiwdr9t2FrMD1NJ31nlGccIJPMaYSh8hj0WhYc8p4H
hEUAHJgi+IPoXjvDAVO9F4hoD8xpoaE6wKSjGhs+nZKMgTVc/7wiS5+C95JhbjvgxonJtiaubA6a
uQaZ0ZI8MudKL5rKYvFskSmBpjwbMhAPsWxJkr+6M8Tm5EQ+Cb//N6puR/jZUukpMzJCJAIPVov8
O2Tu9g1Bjvak2FmYOzDXseNpyEfZqJzVPZ3BLOfIwRomL0xfEhMIPtLgxMxJr0UKhTXmMVH0jTr4
KdGKJ/BhIZvJbl07P3ESlv5WPxr1hIWbpW90NEFxuyvLD0rC/Vd+BCoNDAt9WjZFcGJXPxtt+L7i
E7AEyWAqlgkapG9moAB8itoEqX0ezUHkZFiXpQM7fD5RAG23xkQKVse+9Vgy+CXuG3BUz9Tctz3u
lfPmx4Iz1Ww4uPuGuvmlLCqDPoFgPo09cq6K6E7yPkZpUBCFJmkK7pR7way/LZac86zDRj/ePBeS
sbiUxYh+AoVDkT9QbHS0YLnlmUbHF1Be0j21lon9TJs3qY80YrIoD/geX+rEBPtNTnoGpnvlrb34
uI8AgfPzfudgE+x1CxobZ2MsnXAMO83ytEDtnYYrrLYlVTzZEc5zjPM8uy6tcyD9rxfQowbCOq9k
ldr+eP1qT/0QGDxfZZwJFiST5WyfN/rH4iRKWcQAeoP0heMRV7AQaXQowpLVYU/y0N4EL9ufx+Ym
Wg0RsOr1lz6LCV3fKa22rst6RO1XMVu09if+uEKbfRZKPCJQ+yg6H+O6adh80RG5w3395pt4A1Tt
/21ZXTFvnVuQdJ8Bq/bb/UY2dI3puLIDaaxMc9NGCiiqxo/5z+OnRYHY8y/hkuUDUqO+0YCN0iXw
ZdjfHQr2A2xiHy/oGXpkCmSvFvu0uHltOvcWU00LHpSJ2NRr3ogV+njxHKjf9lxL0QBBLxFKIm+i
WUszIWqw+RUjRv0/v6Ml+5BzSYvxVrAJkiVWDDWiCx/Z0/FDcABqXCqabXzOJiIhmSlVGezGcyx7
MT6VASgwguhStHfWmk7wJdratCuU71D6zXjLUwNZmZUwz45V/OZhsv2LNxHczMZnmfIgFVpQXmaV
0f29d9E4Lh/oVirp2QOMWZfPTq54wHrB1PpJrCWe0SGsL8vz4DaYlx5kOx/MM7vD3Ggojm2OyoH4
HmSZwJajqTmbY7xLXhLlrAY+EQIV+yz+//G1+W9d/ZZCqRTp6nXQKSxnjBcAsRIv4nbuYkbgXgVh
pBPs5SyWxfsGvuaw7TAXEj093KtKDx9mOCWrG+JAShxE+GmAgnNdN3v1QQkQmFrZPONIGzbv1fhQ
OGzd3NDLErdDVnCNKy0r2wrwO4ZFGZvV7HCphp8FwO3DHF2iAZIt2yuZOwMhYhxyGqq6zw5jgytR
mVo0bpzEsO9x1vEbJwMh0OZ4+H39IqnSJILMn/TsvWts5WIfN9PS+3e1FS/I8F97U2gkT6S9/kL4
J3/9TDuCPGMbAj4hKIYSAfZQ3g8odFtB7M6SYBiYrwtvlWT4iP2PnlfaLrPz/NGHTOSUVbZBCrjn
67Z0g80Q+6PpFNn2R+UQR6i7/nb9oTl/q3zZypqBXtCv/Cm+VPyTP5c5kftjlca19QIt5l8MEsgt
QyZUOAfGczZ4yaCdoexxdrFc487iR5bf8BBvYR+9FQCCpv/0ukCZ+GxRk7zg7pchvvuWOaFtwBz9
P/Gy7d/28v4+o/WsSTE3TbTAMtI8MO52L5QjHaIZr/28/UWQdz2oZ1mH8AMD6CQWA3qnHOgNuCT/
H3+ftB9D+fOs7HZGXUWgwLuS3KfKWc9MboClmhnO9A7lV56xrLH42RivlcoAYdImdl2Jyvt1AzEp
uAdC11fN/fRflfv5RE0b/+taFx5rr8YR7mtTLTyxzBZ4vykd74pO6OoWXn1ag0nhc9Z091KbsE23
3MwR7DnXWsF3auLoBMe8v2Fy0+R5NL9lgORtBAspV59LfEdbtAqDmjr0nzaVbr/IU3OyLoGjZkCV
o5LTkMhpVtNh8OK11T2oj9wo527eUt2iiBImi6kz7BH4hwUHrpCW9uXSZnXgebQDtk5Vuu0r8Vl4
vlA1bV4eLaVst51FrSptpm7sTrOSMt0AwphrPdVtL/W6neAMHR1um1nDYWq+Wh9KTT07ck8Sogta
rdHCgfllnAPeFb3QyPFJoKJycv68HyhiC8QeOjFaUI6OImizqRFxM5Yv6/jSkkm/1MtclpzBXMcg
vy5rBDa7mNfpfmpkX163WX5HzVT/cI0ihmQ+0JzE7BFoa0JBaOVxIavlrxbgpYgO5343/nuLkyRs
27uhVoZa7lACoLJ0SjTnlAROOaB1QruKMO8tbUW5keFwWPlxvkn/ueE3okpYslKH4Bbf07AuxFT0
p+HtzCL9ISyAJW3kKNgEQWEJ0wQfM+sr1Cg/2vsjQwWPpNTcPN7CDam7jkhJkT9DII3ThD14oZkr
k1UeNXnv1H7+0Bxd5tNe7vI5getTwXGmEEknkndUn6kbUG07xDb+S+pi6ay9F8YHYQ1frTb+wgKG
m2T7xKadnhTzoDNN9Ofr/gab3mOdnKod4THugYOF9Dx99sjOtNXS7cEf3z6kMFLomn3dRS71Krty
rFzcDvm6r0h/GO5XTG8fAaCVJmgmjsSCj9WYOZQ+FOgHQ3yld2LPDRQL1buzsjtkppb0KnE7ClNS
l9MRfZVTEFsymOMK+b+JvK/qWlObtKDwpUMslAyqNMZrwXimH6RcY/SzDFTS/nRfnSB8Cg/BdA1e
3BYTYOQFseYzRiVHvGPVM+SAbx9uAGLvhtV4MfIYFBigrqE6G+l8pvzom/sHvfXZqRjdrYMs5k0+
2+WYNldI4L+zGwR0gl8Nnkoh5jCb+w5fnomtsMhncZvjOIHs6fHUfweCDgxcXGOd3548pbUNTBpI
32O3q1LzbFD3iW1WRgXtmyGrkj7kH6r5R726JceEYWZqatz7Ma2H79gy9eiFoRfJLaS/LSeNT35e
62swph0/C+ujm9Hbed0qkfJ0aQDOvwQde4ZtHhQJ2G5vSNqScJRgev1adgUuY9gvClfXur2O1UVX
0pUZ19Tfb+l0UB34sT3F6QbhGzfApusMJdvW/F27+qHzerwmw5sh+Q/iCcoxIhp6iEEZK0Vb3jPh
h4eQ+8g9Xgems2K8kuhhjHLCdV+iaEt25+uQJeLfUlRnuKhB3OwzHBshrU+g87Z32OrnC2XNnPjc
QI/04WNP5bLjOPAj59zeh23mzMAqPBtA7tS94YsKlnE0K7fnAOeFrljA7kmQCMBlT8bCMS3E1wzx
+6zn6uc/Gej3lIT6Kr1kJkcE4ImZ9bpQEBt1Hk40KdITxVONpzdrcWa+PfB9SfVBWLw67nHh12zU
e9Ha73ZEW+m80XqeogruDH4dQHDgPf6b7XFtaeXVi/oDKop7Mm+/IBjNIFoR+4uxqbef9f7AOi4f
VL1KYkvQuXbvS2dglazGH97UgerWuTi2v05w6x8ykmv3IUtUqzOc5vHAQnYV4BRwIiDMQb6wBICu
CVRqsw6JLt5TWUSbtsjJ1S6f87Z2aT9P3yfFSq+6EFxNK6NrDli9/eVX+BkwTxaiqKyjVANoIGIP
YbystPHkbciDnjOpQhAZUVj+bfh64rDA+0ltVAg8dDdB/Av6kzY8uq1JGW7mCtW+Jw8bvI2IBidW
WKLdeU+QRTkLay6opaHhGXow7qhgiGgq8zVjZ9KlLpooeS/0Cwxd4u9SHI+qhVAt3Iuxyg83oRC4
mA183DgMsA3Ig7B9hUQQDNJO6CdwtkexkSFjzsznYNPtodwRzQKCpcm0madLv7mQ7sjr8XdM7zHk
b1F2PxmouOwsj4rUEkLfqA+FYSz9UpUohnMjsLDiQUlLnkZBFu/FxRd9nFl8SjrPZgF1MXFdZS8b
g+tRr1mMZvgd2EJO++QILyn8QWd22f9VncvxlFhmQw++xSJCry+MX98UyatxG0ASh5+Arh8nDSKq
lOJ/avvE6qohFmKDBBwZJOTJQFh2wNMUOkIFV9TRRn5D4JjKEiiKLe+2kx9GTNDd00NiCkrNrvn0
l/z24NIE/RwG9PzJHW4WPqtAKfbJcE8Bw3fybCqSLT81lETrE0mAWb15xbEpVffxkhau4UEdlqsr
Wx/SG9WSlxZU4gVPOUHz1W5uAmDSREa0K+pEVOjsKVHWlelq3zCAbKuTlszDVRoDvA+yOKj7DCfi
yeKqJfSZ4DCpop3FRodjApzUbAPaT7iE8KgfcgqIsfawVIWC297tKabPJPxUUXHWD8M+8E18FyZX
t8GGQGYPb+nNpDIYesK2W8QHOmAtmyDSfQZxZRDmljmGRWMpiXJmRqVQ8t8x9fLw8uqGy0u1s96N
dZ2YKqmuk6S/+m1DoZl19o40i+vIs8t5qrUcrJ65SFpoA4G80cWsnIvz3L2Le73bc90S9a7HTWnU
n0NYdOmq+LmRZqjKLmGKT7wUyR+On5I5IO9XgXdO/t9JIPjwk0Vad8diwCjJq+CTR31FWhu7eARz
f7Pe/drWw/8/D9OUvz1QV+599yVXPThT+Uw0wC9OixFTc3fWM4CX+5dzcwGsw2A1vCE1y2yOUOwT
EK1oiN4y0ObKgQxuGLpR0mTuDdesAukUzVqTmIkk/e1wlIt3R2d2oiVpY/Je+kwnIPCwTUA5tkyk
CnjYiddmERR2VqLfESxWSv8msA7Um0V2yUHP7G/ED95rGkaqQP5FgKASm8rK0Uer4XnjUFwEshWm
4bSZpBy6y3YhSp0zT4nCjQvvxPK/FpX4+3mzHkdV8MeA5Pdk9X2qpE5DZZEYWnQs/WSdIfQRZPH4
CjGhGc6rs8Gb2DcQJ6ySb52fFflx4TqjocAErhNkP405WGFSwmhS73ZwikRoZQN/On+/8sh+RJp2
jP5LPFr9A3RqTsC1/FMkrElN7qDbv4CBQikDZfme4wFiBUiCPmkqGDxEoxxwe6aZbEIFrFdOxJt4
dQkmixiFEQzIgrXZU/loWa75Hmmk6LKy3z6om+OOOvbjWtkzD94siQ0euLmP9ZR7GNf2ruLgW+/j
GluIZqROtUvao+yZtSnaIKqq3I74o5sZ7DOskbljDY8EmAJARaEb+96Sc7/Cph20xZT5uSWkq+4R
r4kGuV/qOjT9dkxcydyqDe6i71c06kPC3tAhGJdI4qgF2VPmKyd6zmqNTd1KZbkMBCTTtIV8RIkT
Jbc4JYuPJHfKYhK9v2WcPOZgEoLvtAUQwAmgjaXwH+7fwDv34nyZSvlPhpCWIsNgpIMeak/CRZeq
rWwAfcrTgpOeE5T8ppRq+hRzcChaitI+s6gzq1jUKHahGiDBSWz2mbNsNCV4WUtE349f3NUMQbsq
4RGut2hPKYqLTL+dZ768urXyN9geY4FiSU6vQ9atFkE/PZv8Gc+mTqiBuUobQByAycVbJUiG7uVF
h0FY99OWIKPn9HkALqQWQxIVW60sqMqSFyBhE3rpJaGfIIsXLwQunV1VuqRTj7VueMWFifnezv2I
uSuxEDY+RJgftDHF6nQTO2FPT6Kt54JQIWjPTHMu97T+e6FaMeEZB+ubwl4Zo698V6T2FSLAmotP
KoU5Rs5tBoHDIGDHz3uPIWpMUP7/xPvXWrOPR6+evgz1Uso0ePIHsZDQXX8WzAj6tr9kg7fFbCn9
1UOrUgVCYa1Ee+cUK/eFwaddXnLhI8IDyjIADWCRsUtFfTA+ryoZzajtIc9r/ByubW77XCCt617B
6aHJNfjKYAh9XmVAM3OJ+ySRz7PZMTatIvhi6Ta+GjUtF76iM6LLEe8oeLDgYh1ylNtm+/RtVzwJ
jZjMC0RFwoczzcl985kOCZ19ZwCTQYUySvRq2TFWKyHagC8fyspH7UsU833gtsLk4iHqitWnXkze
ldDTFYsM1tR3aR5c9WQ2Qz9qoDtHYjfmcJnurlGAvnNM12XLRbOChLJVKNki0nGEaa7q6Ze/nsLs
ONRDQGj85Tfj/am6h8fVaTwDc40y0tAB0JpmBFhxxh4igQwrynL9gxESAkLV+3S0Klfykq5uR3an
LzpaJurtd1oOPbNkCwr2iZmbPKATr1J6NMcKYoUBKSaRxBpwax+QE27Okl62hZgP8bp1pfbJxXH7
bpanqiRwG91sWrqO2tW6Y0E0LUtxyrGZWKiuCrZd1ivwSD2VGfdIuX/mTChycnBgY3RQxn+JfM+5
IGD5w0bGXnYw44bgue4OJdxrmZjrpN6fbRYA6VV9gQh74IEh+IhQhd/Nr6NV3pxUSp0kKmBIehwW
8I7unP5IYwDYp4170OrEpVbL8CROHq7Ldyz+zo3J35Zqs/OgJAGRKbV1dAhLIJ3HXcn6hpAGWzcG
ARGlwF1UmdptF4NVMiX30ES3pyc4fH2G5h700fooXNM8uLpVKlu316PPC/hlxxNlYLtnNpS6xG2D
YvFISVNUNc/jjFyDgo5dETsLPrQYzlVeSpFa5jI4F4wY0PrUVFY38M9imZRyKe5NzQFvmMP+F0A/
k1Qgg8kvzc0MF+iOkCCC1rODW/tzRRvxK6VhNUYPxSKDeURssyOFp7EYN5iHGy9y36QDz1UFo3S7
rO6oYEECqvwX60uCMLkm2nQo2ae+21mnFGhNSxYHymors2h/Wj+Nq/TYSyhvpLOECSjXbmPY185j
PWJ6xWk1wvXMMqo8cEiqF44cxKHYARDfcPBal6r67xlr0XmL/QycsYt5/iwkJidKaKImBWl8+9LD
I6fRDHPoq23lHtItp1zMQ/8pdAokrTf8jgBqk0558Dw84kIysrLRLVH42haW0nRKGKK738Zke4/J
IZY8sSnKROiqyTvWMu5dWPRmcvNWUinIrFwKsgemwqvpxnEzZUnnldAEhTiu7you0HKjt15C7vwG
KGU1RPhi7l1IkOMe0uXjIy4Jpoa6++wUMot8tV4TjZlrCT0tDDpUiyM9A9N6dj4lfxVEmE/MEOx2
0AfuyivZDKLkqyrpgqIms2tt/PpJYnD3rj31xzV9RvxZJU+5B7cf0KU0CuQALE3QSJ4sa5ZxUMzZ
+gwBD3mgTnOlXHmvVUv1eWO4hLM6jjaa0JChy6xEa2EXNqljL6kYKzc/W1wUwrUY8EUx//3V0jo2
oHD1KO8tD161zftoF4ErzbOoX+/LOBU9A0NQp/HBavOg/B+v1KH/196zjOtBttIpK2O6wjQDlJf6
PnMH2gZLDMF5KxnNFnr3FcyIKxqPaocvlGJuodFof+tvL0lLwSM1B5BAq3ZxzOS1vgnPUxK7eC/d
cACJH7N3D/JFheyVTaFesbdZFBZo6hsy3UtfIbZQ+Y3TlW6EwShJc+aa7EAsBMQLff+67LOOXFzB
B4eVAqNuDPLJZktRNkehGT6XHEtFZI52gZOJYhP90tdWnLTo1jLkcbK3cjk4kw2EGcMifYxjpuyB
vCCqX9WoyfN8UNAbgRedRnDPsWffVqZomonC2pwcoJpurueLpZ13tb5bWN/CsuqTX67t/INOhuB3
18slYhihreHhd6eOMHy9d9yFP6w9yS+rIdVENTZxWune8L/dcsBV4oY5SX7ABANwsKKvY+5oy/as
P4ocBeDdAQyh7My6DMF2oes1wiYlFa2F0YgNAftANLIBXxvr3DqmkQCgscOJzntCAme7QHAdlAmC
2BjD0w5LSrajj7+qy5fYFpoqAq6XqCu0HaTxz9ILQ2NEI5I42pDXhu7q/mVGEi0iywOKCJ3lPKyg
3ZGo5jaUd4q3bL7MzjHej+E0FcwjbeU2XhVu7GkA18YOvvPiwsysEQKKsC9/KpFoh8pUX9q/O6WZ
RzJY2qr94hZG9NFYdiW/sZJGOHfgMUQNBcgkG9RL/665py0HwZEZv47ZNl4ZyE4LraP5bG2iT76X
NDHLiK0GtHIQkIPTnBN85bMmVEgyFe4TnSegO5VjnrLqPtJUlhd4nzAdEQO5C2kf92MMfZAIoBW9
4+VaV8sDbGlUW8sC60eQp/pwTx9y9O4rhAp6WHKy1SLxJxj6S0T9OOYGcuCltY53fnVxTqtokRif
6YSL+PnH00QTNghaXndAJXwIVBHTggHgqQ74RsLBirvMuY/a9zSkIsVB8oxFMw4B+X9MzDYNTCaK
tZ/jq/ITClh3T6LHZ16bEALd25BmRM7+T2OT/QBZx9GhmoWcPvnXocnbn0V/zWrlcGBcxS0UIiuo
AOc31yYxNW/L2MOhCH7n5C6zUUIAwUcUBxEidMXM4czokcy/s8BClcKT516rafpyN61CqnSB54zi
nG8DoHvjGvohpaeJ76OwlHXeaYOqNzpTbBEemKaDJIpkXxCvjDqQDiX34JFD0S77Aqdri/7ESAXM
eA2QexEFZwhFm/nKgNRXRSoScKNbLx9K8khGJX31CUy3HZ4YgUENvkZN0Z9B/NzGVuvF7oRif9pd
MRPZ53oYcKa8GDBvfSDx+Tf+dbIxFfFBjrhXHnmvD0O5PtoR8vpzA09vXMBCBQulqAkkZmx/jHs9
gP2MxQv33r3DkS8yPU2SZgx8kDC37BfOTGLffGOKhu+YkPmg1DUChDsCyMgBYfNG32JrCFhaxT17
fbClk5zPM5u0qII807jjVsvPA82Lc7igsHb1P70l6CtUajWm54XXqIZbXgpRkKVUe/oLu2OaT4gX
me1svffHAJxTGNOsIPzr+m9dLSbYJ7+zzrw/oQrwb+oHXmrHPreQN+G2LOVOAhtdJt9i80aM4zRT
UXIWPpumz9oZ2+IShbEvWfU7WicKIB3idY+4VnuzS7pg/4TgMhdb0d903CDc3U+5INn6DOV1t6VM
wcZFPEbhYH2435mfYK+T9OvEUSZDRSN9PsHK3M0/o8qi4Z3oZAtWMJr8QmWYEXDUOjmE+tc4vw+i
cExa6cFMCpwqLuKuWDYMfPXx3yAh4IOhUFDj2SkKEiMIi40oiAc5RFiK6mRApF2il94SSBWoo9bv
XK8AmLCxu3SzgN3Lqi3TJrQHF6U1J9QiiKAA+i5MdGo64/RmlwBfkhL0Q/vE6lGpTS36SoxKfw8D
KXpyyMHLwuK9mLiwrlJz4kG3FsGXzSGChwmqj+Nr/eu88NAKL44nWBUZl9/cMk8wDzfaE2x//Uvd
1E698rU3YcFLbdnOuqkjObf7ijXMigPg4yBD3S15k9YfHnYUxhOfcufCAXliBQ2fL51DdgGyBrFY
AtrEjwDg+D+7FIMoVot4cq3Hc+Qly1/h7aVUiZ1QBAotbJIL8q61VuwGOT5ZjSFWqRyXT6wnjaAd
RlrBfHGHyG/tWYTQ6+ubwapAkZuZYzhnl88x7HZTGMSG7+bvXfX4mF2LXwKV1QgztvpyqCmuDQMn
U5UUoyp/Hlq4+DuYL1OX0HyGkHG43Wdxx0gxVQNmsrVguUEYNh7RvEX2E/02LJBnmX3EHP0upAmk
om2BAE3BjS4sXa1IaAqvvkt+pE2yajwDPrKKosU6rft4WBmhldWDh27aYlnf9A+00lLtv1wxPyLU
k4OBz+BGmUxB/qNZHCL+a5PI23qZ93um9kKh34+BUoVkV4m7PeOxzh+RcTFms3fPbca5ETrAmCDj
v5WyGp1zfFbLrQv+d/KfAnY0KxN/+X+WXoBb1b8ydPuZBJAfeq8TvUQ8AzJ9glUZ65vdAv06xUAP
zwJdEzEsV/SXZF7cgJ/moicHjyzKGAoXs5JyAIVOyN3WzTLfA9Qu8Fczvd5tIYcb49UrT/IIPJ/L
WyolSa9RzXDjw7/Zjn/wSwc6pIRkX/BXONXWhMtugKffEokar0s1JK34FHz1Eh+cf+KdaPtsbpy2
opGR8kEezLnebHM8DqbOtfcn7mXaHgqr7i1BU9qND9NZz/b4oX33amjAKQEomLvpmfyeOwLk5gGo
PwZy3V9phxs3y+ulYRtt/D9GSs/fVOXSxxN4a+ifARr/cPp7ANOL2i1hbJJCA1d8rgJTWEVR5GvT
0XVWry5HKG/DbZywSGqSpXxl6OxnHIstdjj8ZMpOY99WpeyD63i76BBq/wtO3IybIdaBAtx6pCKR
LwSKhaRKxK7CpynVsdaB52oRWXR9h0Jjgvau4WepElcJhq78cKBA0twdXvH3xIptrWZWDfsenLlM
IdARjEdoimpTWvuleUu2x91A8MdjIdcla847+64sKuMRLW21sCYQXTla2yQZL18CYdRhVuyI+D1h
jcmcCHyD+DIc/gw4sHEnAomiVs0oY7P8FlTsBAFEq0fkuhWbqxdDAiyNL/mjdhcTUO7enPX9aZ2y
0MhTlfnQ3/pkp0QzDmvvbc4C46yi1BBTzfmaM3TBc72Y3cpl8CN4rjzfIqTQ1D85T9ovfSslJy6C
Ck/KMw3hqYaiKOJ5LqLjn7oyzg3nS/zNwHS/KZ3wmrrs7NuMaChUvMCIRIx9V+CK214dg7qa/OvK
jj/nP4gQK+viYMH4Ci8LmL3QSa+dACugv5Kjj1zq8o+xrEJTsq2Z+JYwxprsNBu2HHXs1EXL3Ffs
i4srawwDUszYGsOoHf/hwBD4HUSEa0U6EOldnyf5CVQ3vLFrcCyI/AUCWNKHHjIvq9F3RPeKUsS4
kYlCar66aYiY1LluQdM6wBdfGNmE+1aWu52Z4pX1qBujnaTFECy+LR6mOp8M/L+SOHQffEwf/QG0
UNSK4l/svpSY3gQpwTb06stdhD5oQJzA/ZrsUzbFAan4X5UFM1tQqL8tsWHiS4C5/q6uzQGy5oqs
YeUrMB0OQX89OOFMVUW05fEWaEwrtGw6BqwqXPRAOwEPl8U4ywiRX7nKiksXQh2GMhhWUBQ3kR8D
pOIbpSbGDSewUdcPLDpxa4Qbq8r/zCqA3IBTgeIYh3Lfh9TdGU8BKCy5qBadDLBkcffQ4IbobrCS
sDkN+x2KIeWKkaNXGF0ufNKDdyFCSnKIchJSvAfr7e4Y4jnMI2gIanll+OULkWcqmlevo32uesbb
rX+4FjPq+DkT/mfl9KTHC+j8zUUkmKjUwkFx+8fUeUElnPfqh1/3tH1sM248Wa0QtgtHU0gMPlxj
imzFKJhxvjLH9VkQr690HVGeHxw/ExYUE+9FHIKHCjDHwolFAWlMjx6Gg0FJRmLDkOwckd+DVyKF
9TG/lOvWbCyXEL4VmqrBZWXCwHm/szCii9/vRiRKTywB1Skt+pAL01yf1MMcJRJ4EHP043amWJPG
Z3p9YrP6qk9/LGrzGq93TaXA4oh7iAyVZXldooiyTrBbQZw1yVj0GQOg7NCj4ZiON3GCtTS5pdVA
dFe+e031j2EoxulyYIFmxXkbgJUyIxqFY5N+Gj0i+BcbXoLXGvmberpQOGUeEk51TM27wqsIVpXp
YxWRQIocJgeG32uOfOC0hxSViH5SSjMBkAMX+lvT/9SP9Uze+jKS0f6Ck0GcZpDpo1736awkZ5Au
bX5Q7tKWwqV1nIbtu9hcTR4oKqFTHxzzQaS5Aa1evxcwfqLwHv2eEd+O4ivwDnFOfKV9wgCZY0H+
Qd/KtJZA33Jbho8m9d3pAHroRmFb49iDPSR0CoEQZFu+NZIUY1UCfEGR14f6X6mw+xyee/D7rodK
kjLdXmVpmflebLN5kIn1+kHI2mM7y8A9f7J23A42pLtoGTmIPAHYO6JI1A3bKUsZsQuT23CU7YLr
xisqGaK4xcNCLI8WergZKuXejCLxBdzY8avUtvaEGsdRLBA7dNeZmQhCMaD/tf/C4nLLyLTClPNy
8J9jQ0oarJU+gsdIhFZ9+Z3UgV2gJDgwT9y5P8x+W/Jd4rz9FEerKIz7pJwhFIUH6sbxDVcV+dyr
K53XjMVZzTB4Ap2dfw/hKFwdfq8K01BwbU5K0mgH+58E0HBNoKQ4w3672E0+KbIz+VpOWK4F+N1B
Q0DteUxTIDEdu1MNB8bPy3dWFFiH+ALMf7Xb/NevuYEH9QgXdjJQwt1aEotaxCmDw41VntbwZ0JZ
ypbhFU9mf/SV4Vzfduz2vaGfN79Lt5sLClcpyAR84EiV2UpiVIG7pF6UcNBUoF6MngTDGH2Qs57r
3upS8l/tV+d6dtB5AyQA/79VQPAS74bNS+31nncdCADuYWLl32Io9jh88EgAROT61GjJasehUjR5
6mZQoO3mfvcvMf2CuwzsoFYMS+ILsSeETwqa2SUhCYVgdnNdEPg/aDgiiO1SIAw0luKVKZYmavyx
WJbeiH2myx04fyS2ePQ2fmETXhi5RneULK9JYLMocDH5m0DeRDGRS2q7MlF/492hwJkeM0cXCdmU
9oFD410IMiDCszsaeyw5MyFK1IGGzJ0MLIZlHUzFhoeDWVj5JNhA53uPLk9zDK2boA36q9b4NNm7
mdQkwg1bg/6pZTmfcXQZgXO+R+KwDc/nhGy8YiKmE1sHFZk82BQugOhDqBMHu/T+FKD8i9ThQqWL
kWLFtY0Cuk652BtB+wt6tcPS41BDenu5jYcaXxCH3vucES5iSiamKl5o+7iDRlZ4DLuT2PqlaH1y
Obsri59EFq9Q0YPx9zBShFEl2Yf+z0vI1rnHJqmBIabNr5kdIP4SiKy6YhdFz3+2WDIU+JLHYnp3
G2O+AK1HZh7OpRLuDHNQz08lH+gTIyCEb9lB1FZEaWTVbGk+OU+/DyoTNgGEAwCGu1rhqZcRfIL4
ipLZ5WiAfooXKO0FLB3Hso5R6pirZyvO3bPvYgcdjoA19PHdvB2/kIpW5vop/Ld9gX0vSkoodNfw
xPobxm09RCHnkWF5aJRbh7P/rG96mhlk+trSmUKwHXCxTqK9oMnUhDCLlqq92LbtfgK/0LAqBwgm
O0rYOQgWWPH2FyN1DvezcNcW4Ws3CDVKiXezc09Y2Hj6sKesklnZBhUhITl69SpUojJkBmxZzlpt
yd7IvAGgc9MYi5wYgvXeucJp2bAvT+5QlB5k/kx3RfydY3qEm2WgIG45EBFOU0nJZsaXoZLCeoA0
8bPmg9zfS9fTse2FfSFqiKwGB+7B7ozVTG6A0QvaoQD628oXGG+ROQhGrNX5h3eizRBrsDBhLurB
sbJHJI7d7jJowgiTyzIQkFU72yRCaRyHG8b/wgjU+2pnFp5InWut09ffCbd6na3oblGfUwrzFsDl
/TzhxUUrHeri6M1DbldkC0vQBHwdRlbYg3bhRL4PheOIZfx3qnpdqrFPW/QtSEkhp+Il3Bhp6NH4
DUj3M6JZy2DU+78mMSb7+q5mp3PWbtotmgC/SMrWn8fx6bKa2ilMQHn5k8O9/9In4JjgPjSM5UF7
PkBSygBqYS6VhX6o4L24aiIsYU4XZiiBvbY1N7VWEp0+RI0PTPM/mDxLrzX5SqmHJTIR1OBT5T5c
RB1GSofsLSZ1WWx4kFamTSNHXNudwkAdtz7HQY5twSkliMurYI6NZ+WmsF8lZu/59IlaJJkXv83g
vUtifKls9p/LblebarSQnoyCheJ6Ek6gDBNu4JOnhe0d+t77qShd1h0KrtipI9r+j+OSZoGJ5v4C
t84RayqGd8ZLL+NFIjCjXDJjI6cCEKq5JLwsswWEow4AwaXtIlMvYd0tBGqpNwQa2AmetFKktEZQ
s6YiHp+rlJUNzHc66uHPQ/HjszA/zQ3ZsvOWePWKdOTK6mxyTuXWoBJsw+KY0kI5XaYC0QykRTx3
+Cf1vQGzPkFS9PrBco1CJRZ62Qc4lPkhzDgdQbJhGJAd38kBXPHTbyfP8zN2vuoo101woAfzyu+H
c3G/cxlPHEe2UEEaozJ5r/F3aIHY+2/1v32/hNeWHvlYlR2iStm47ShWA9vxVHB7g77sbO7F+oWv
79wQ2HuUh4o61Sy+N976GB9lAQO304c4SGgowsuMGXrQyA8l6hUYtq8OEgtmfYabuADJV295JgT3
l1R8sqKeRFQpbW0z+e7H7WDJIoU4INyla8EnqokSI+Sw7mMDK+XwX8Fs+GrXQHH0smz/zCm3xo1v
+xDBylL+tCHT4DPAn7SVGxbfAh8jnXlY90fJp+rdFNmPpnnktZ8UUJY0PAiJO3yqnTr2M/uPCpdG
U5vc7yGq6TRDJQCmE2ZEkJPSGCdDRW8ud77jT3wVbSD8VcJEJapVLrQ+L0aLd/TJlO9s3meTb+ii
Dkbex5tyDiaAitg51KtyUOpQRiuLoKN8LBggOZ6XP1nEM2lKfjuJxx4S+YReUjhzPUOfbFXZBzKQ
dZSQqCKnjXZxMf3uCU+OGfLYajdbxz38c51E9LZjWHtQpSw1E1m2FGz3iChxenVo3b03tZOMnaNV
pNYh8FE4UUvrSSZhpx2eVJG3yLQLjiXWt0zRilTxRLLgnL8wPxTMOGgZaxvac7zTFc6ndDyXopRf
PTRslR95sTPj6q1vMw7Lk3gkPno24I1yNGk8XfOJN1Yj20qRvc1XxaLz5W504P1fe8haIWQPi+NY
+yZlwXzBSAA0/xHKA0JYTSGhYU0nW1qAknAfTs6WLs3Lcp9mC58tK3nL6e42n4dP7Jo5JktgVSef
gQDHdaMJ+oWk0+NKLMtVuA3f7Nq1TzckO9a+YLD81zwLL/jlRRpbkcCcsZg2Y3xV08c+5q0PL+6y
Uy6fVl6wITFJFA2SKWQMNSKCUR4G7SSE1ooD+2hA9/A0XLwUv2MfYOqPMdfp5LnQFfdHOQPgwGdv
pc0AZuiU/f62+pCFajbegf6lQqv1xNatsGs1uw8fdlyVic6+7mz6mD4FhbH/44Wi7TuFRPpKPY/r
pi/enHPnFih7ZQ5VywaTPwJEZm+oFaTVifXF4OiWuiYlOw+zI5pUHGqowUgGgJT4l4br2m/Yjegk
aSALzxgZCbrCthtLgWArcY1Ii9QStZBwMBCiZVviIO/C166TQwCGbOFCjF5qsOubK8iB8K4USaJO
yAPgg2QaOK+1siQ6r2MDy12IJ/vIHEX+OwHN6N0MeOD4CN9fqvY/Itg/IbyX2q99y3dC43jsmgvE
6ySr7ACLkP4k2asM1RJfky4jMy/FUu779glLAa44ksCoNrbHEzXgebbOeMXeJ4Zxsq09BRjECq4c
GLVuQGwDtiKIH1IAkbuD8WVCzHlgkzG9R6FoYvJShIBUxDJredWm7mEQuFUVDpujIOs2I/Ze7rsL
6aV2o5rDVd5n6dn9OInkufl2x7+aQfzRmbY5tJM9pugxABToybHF7gjYt4xH3fM1Xk0nQpaaSNh2
vfzlnt9wSMcYkP7arDhZsXjTXnnarhy5DH7tz2ztNEq0ktSa96pcoljEBqFJqnW7AAuX5bNRgqO6
/kyyhK25tU41qkUN4U7rUimOGVP29TvXkfeLJuOXC51HnUK5zRy4k33q6zvQTexNmZ+uy03IRPL8
0YmDM95XS0jEeCMUJBsdxk1j29ChwRmdsSq//NF1PylmTn+vrkn5MMALIkSNsf8iOJItKdZvrysk
qlXo3aRGAvf9EGf/SNetI8gbC00bpJX2M68wjDD8Ee/NdmnXKYNkx+ZHkgUeQuHbnQG9sNME6nX/
8jI4dQoVZ/65HWrNshNX6IIAYycM3EF73rRkGRmIXrneZ6FLf9gvyBzuJqRWkbVEVPONjz7SPpJj
VTxn73ZZ+dV4dlKzQ8jHgWID0zcyVqrp6FtPfoGYHzvv5o/rV3Qx1sldIgbVTwxRJaKovFkiEULR
WZoXCUcheEmSWTJc717sxktZg2+Wh6k1OzEab7+vGSD/hnHeE+oe69gcFuSvIPNT0AUJpxe1POtY
n3cl1TeVy5hH/Z9m5vAbWLAtZkgnxbKG1jeimivSgc+MmRM7QGPFaW7pJ51eTZpt0xyUY63ghS48
1NHhWGvuG3B35axCY9orHVBNM3WnhzEnmPuKlWW1ARfE+KA80er+5tGu3a2tvqGB6vkSV0rrrSgX
01n94FPj9J2sNthYz4IoyDAaaFtHR328XhGtd9hG318BBec7KLz3K6wlP/8nJVzYc7HEI66N90ba
x70AEHjYuAJlHz42xKN/k9W2vGKdhI5cgjMe8vbtaCu6ngfQljD1zRnlvVFP4TAZiUVC1SB+c7P8
KorVDZROqKHjKLcEIsDLTCPBoRQGQ4q3lazFJY7M/+PwC2zf6Ih/WfLsYEV4jMECxu7r5CP815wr
85lQfWyJztA7Y8TtyTb8AkCT3FU6P6pKV40F24R5I6SX+K/Hp3BRys312cl2+FfhfC2WDy9ksuy0
50S0Eq9CU9rTI/SgHK8dqT3OXlVsvLzfNb1jF5ezUq3Ry9nrz5HLngWqvJ53gmyRQSmv+yuNPSmy
SKTzrTE2F97hxwEwDrPRPs10GxmkOsqHRll4oYJKtudfIm2T7eYdN61YM2ERy25HjoTDHp82/p2L
XWsLpyu/jlpISTfI+X7n2X/FUoqfhok2JchepcAuMGgT4V4XZp+pApnGPPHSBFs9Z94UhOL258HI
B8dB3xKiDZHuaf4bQzVbwLo2oPGQLAnpwVBHhFi3OkqB1cAYfG66J0SPQxKBqicUMnOoHylwmK6a
cmn+nsrTkGKIIji1ixPJ7AcRPC4yzSQ6OFiryuhyoQZy43gIUHoIG7b6FbTgsaTZpHuODYZN8BTY
J6yCFo2aKQFSmobVtuTOFN/a4ZXVAPfdaoI2VzVDNIL0AyeNXDQnqH+DjrHjUBT4fS/lj9JgjocJ
eF90wPxqyimE1FkCIkqLZpK+9qVZeWKtu9r7xWrAXp8CgLNrXyHFfO7zGcx9wgkTOuBkE8uoMii4
6ahzNXk58IWsq2yhnqFicgtdlP6Heto8z/Rr5Qyhn4RjjL4zDH2RJV6YMISFJNT8I3Fac9Ki/phx
405Ko7tUW7trIy48gUrMoKl9zeqFMyuAqWmhN+PEGhze4oV3OD9+DY6MdZCeTdbJATmxjLfk3KRe
xecZGsMQ06r+Br1cAWFx6wT95+Wiuj6rZPX5L5mb8SPStEWyErqwYG/4Z+ULM4RjHAT3MlVKPPAp
AFZ3Lw07Wm/P1M9l+ZsrqvU3DPhiWhBKHGR8kE3crJadqNFZbsTGVkQOfwg1OeerChv92PXWN9gx
tObRqgWhyfXglJ2S3JQ+NtargI5Ad3WPP3hhGurr57pFZMZM8Psg3d9ilYIEZ48ikqmnvtiG5puG
2AK4wfMyaTVQbDROJk5stEsZNTuZqDebLNc9qwZ5upk5T00pLiU797Z1hYOTsH7pEkz+molXHvlG
PZb3jzMZoHxG68YtLQ11bUvsN10XzGJHo6w91zs0MvpWdmk4UJpc6fvMGkrMEaPyF3VphZ3GPCwz
PpdLz9+HcqJWQn+DMt0+8aPj6BDyFRWHWd2Io4Uv/Y3Vb/A7AZdoDfWBeaicemeZdCjcfQXdoCVI
KDir86dA09apmJNj2n0izpDzxlg0M5cp1PSYfvQCSIoYk8uotSaI7G388XMLh3mLMCZkUpA6Zthp
bxZjIA63UXlhUBlxNjftVdxxK3UWTb4wGY9mYpcR4jlXawgyJL7grVUDHfN1zX5vpTiL8ixdZcjM
opo7xljivcr+veqG+ET6+Uwt+24c3Im7YeFnr3S5oXj7t+X5i6gkhtNclMjEpLbpFiWX2BQiHZHv
z3WSux/bGUYLB2E0Mmn9S06ahnXfoja6Ehw2R9cJTN5FOkbDEnIHP/qOjx7Ij6BUwLvC/669W6ie
RaZND85c9xWMbP944f/MdnhQdGQmzZO0Bp/h/Vi6gH9WckZrjfHto6Q2s15cResIuObK0dVU/LTY
Tk+SmmyydUjOndE9HJeFATmXGC0YIV/+JoDTgFjP7RdPFczk0E8GLdMVbLH5+J9QcFvQbv7wzLju
D4/mLl2S55kGT8d9k4bsbOvH8FeZVlESaDRtOyAXCjV9MeThae3ZsjD3xpEiBr8OhJwZrYPA9zKo
T0T1Rlzo1/6lAvPM8mnihRbog1bSivjUlLTgBJ96zlOM8ckdXEml/vGw3uj8xz5FEjoIRbXm2jXy
ZPhWLXnppm9mfHRx4O0/bOhsal3jmTO8XpXuSaX96JbQSNbfcKkmwRwG8af09bvn/4Mff6pCwMhK
V0p4yEYLQ3V5Z22PQF3E1WCZDFWyz+TnWF1lFUFR02cMqf3zP0rE5W/J7DAQLth5ZIdekox6tK82
Ro2oKdKQ1DpiydhWwColAPEE/gUkx82Xturjz11TYRxAWvbsKosc51f4ahKtr5h2KyX0LR5NX3xT
NHmUNm6JWEAsS6qGZQa7ot0Dle9blmfHuqGJtLQXYCuYMCj4AlXCWF2TUYivT4ukyJiBfKM1mGbC
9lgukk1EYHpcsaPK8/IG8KhiZgmleA35qFoN9IbE2CHzQt9tFhAKvEiNuQYxd6mFRERu+j9nHt2m
t3HlDPVQc3poW49MIsDcB109qN0gN16z6xE9/UdfiyySGGY7X0EsrFe6vKnBF8ofEZRmFoZIKc+6
+NMKZQdovUT1DPQ3ztr6vEBNV0grBOMrfBGuMmdy8WdCTzOvvfaQ0acOTv90qd6Rqkf6UFO8ytA7
XWQkchYAowOXTStFrRfLVRlMNzn1/IDfVOGaE0MzrF80p2ovMuUzfrQq5YzxXq12UBF8ZlzTbnq0
ArU2GdLZoOAap/5/AXABHU4AmHrP1nuNWuJOLTsn6qBa28Suooy9D+22ptZVPzMTORsRg6xkhTg/
jgeS+nJcheKTv3LTS/HjiHy8SLThrJdagPBRkofkPmS1sbiWe2uVp3QMrAou2XjrvfAJZFkTQ8Ez
J+U+bGRW8q4OajKpFQO6Ly3mQVxobooHUJPv3VCdDTtt9L7hvpkRxzWRppKyGtnKP2WGvaQlYTiY
YvuFXmcjAc0/tUNMC99wdboOCsWec8p1bDk5B2OQD0GbQcuy7pSTB0BPNoKjhVz8MB+9A3rm/Kmf
XbXtcw68aITsCiIWMiVoWTrmfacXx5M9vqnEDiYQmBtQiIWP+m0i7p5dm6JH5OzXWvGBIo0dcmzj
OMsWQ9R+ckUS+jMTDVQ8IIojOCp8E9i2yqUMIibsLS+EhSmMbHQGvwqzwdKwCNRojMYsAmqVd3X6
qUZoGbPgOIRKALMJupoodp3OSM6FiUDea2Cz/d7VRrckkJKnf9Fjhp7NKmXm+NpPMm0yMEdOjDZt
t1510pvGFs+f1gX1uDVBMygiBn41wuoRxhF4cDcp/smxchu1wBqsxLaLHz/+CNuX1n7O98ZJ63Hb
6qj22OHAHVL4IXpv5ONG975+a5U9q3S2+NqP2Q1C9ofVOFyU5y9Flc/PbU28Gfk1b05c44JA7zaV
H2d1+k7TI3FEuImePyu+dSDEvEgl3dtQqk8xaZkBT2O2VuROBbf4HAfscbmTB8jK2l1erDS99Jgz
5XZ86k29OV8faa82ZWOpLrr6/H41K04yIBNchCUDLMhEQecAtblOoj7fvQuzrdHekFDXqJl5cemU
/Vgh9i4q15nRjg5tNugat1cz+DMi+pp1NhPkYQUKLiq7xc0gGJ85vGZXDpAcvNQLORKp3T6GJNSV
/R1GeDd4U9PHRCrdB+sC0MOrJ/NT9JxiTFSgEJDwul9C2ghOq8AbGdt/ctW9I8sxsLLcYMsu0/rM
5oo8ocYAV0J18HibdPVk3BN0lqrhGc3EOolCBOfk+z/5X7FliQoJxdpII8UeMzSk+6W5zDgwOxoc
Oso+g8CCPJsFgiJy4LVZWJYGP5z7tbRdTi2KIYZ00WZOnirxIauZTT8a1kFf4kluzq232PH14HYP
mx69JAmElxBOSVWWLtA/Oz3jH8bg3BueyPmO4cJgA1CpM/OzKJyEILuG8QKFzok3jH2WIIrJvUo2
LbkPBc83UvTm9EMLSw8S4tUrP1ERTtVfWtENekH3P1u8X017sGeWIWCAt39v0wyD8Xw1XOnA/b/n
mxJA/0M1/D+BvbLAnMn8mmz/sqR8E6RSdQeE3vPOevaRMqshw1HQclEQ8LF4+nBXb4ElPwZtPSAv
jETfxHMPEYDttXGzqEDqJzfF2Cwj1G+84yJvLaswGh+dFSQV2ffyZcgdu4XDVIC71em5QyRjBcdg
vrurHDsrBccqWZFdRzOoKEeYtuXI4jRxmqi+8qZQDni23xaXUTeYSdWH1E5eJ2RnNCB2Pmkm3Zom
JIyGhPS/xiDM3aTiFVCeQMn7EtMbxV4RFwPTxdVBaBV05lQ8nGIOJJyQXHX8X8McE6wSACuCu7fM
18bjTStQQ5xuOyM1bp848Fd4OliWfWspHLOmFQlDZYZSHzdRrxCDHXXNFN+G3MeA0s7W0wQkIdl0
g2adrtiSoonKxOBWl3FsyKOLcymwbMXJD4OV6iNQUiHkZER8K1Uxgx7axQ10ntjmeCNnSc83g8oN
hl82xNF0432SOJJgIaTYN73yAV2SosQG9m5SNWcY4b17dop8lvEe7JKbhRT9NQNRj6xgXvDiDCWW
cgXh57r+jnjZE9AViXIpqY9XRNYZDeCrJcEYEorvGXcadxocSq9+SCttQX7JZRrsHBur4U5MB+ko
6b9oVOapN9EwsT0woDlV8qrtSaKsAxzCSDoIErgGAceF2yLv/7S2tY+OyGayg3dMRqkhK66dH98n
Y5OJ2BmLScmb7GoMSpPrQSM+x10Xn8k5StaOIFvHyepVpfgKJoAUpKQJ4y10Qs/Q7/I9KjEeXptW
mprqIGtxdBqXSB9NjzZR1YCSIOn93DQEFDvLoOUDc9mPSSnu7/EKbXdnTQ8mReZQIAFZI7Z8Ohmo
o2hwyt2bhPbNweWFGWBuV0c97UfZZH+wJu17fhziqt7rdzXdKtzCUn8HVBwjmN6ie+gP5ERIPrVy
AAFZROxLxhLfLvfHUveE5u31YDyIeatuLLAIdKtugPc8SwQRdoh05tL+0DcA9J+EDoMD38o9coWZ
2Hm3QB8lXm9/kPnezrtCAE9/mF6iRZaiQMRxrS7AQWRCsaBkgHgXtV/BSfGyZmBe+QMPFX3By8l5
Ggn1g6L9tW3Mf4OseS535cIwhr7x4i6muJgRBYAT4opnmcLXP1UazUL0sr671s+y02Za6h7hrJPR
cHESq6LRGiTVPNxT9wgu8MznZ6okeLkrsfB3LFBNfagWPfFR+OP+xPJd6n2pYXOm1nk1qZd3chBa
yHhK+Fb7jr2ObPb6cvbksLndhLHfMWj+aX54xM2n2VQ/iHEvlC1HLvGv2sLNHigEF/NF1NtliTo5
BmPga7RHjCoQBlnsZONPPpCQ7LV3DG7KZU3baL3eq0R9K4rgQb+C4jflhp2BJGrzDB6GLyOIlDCI
eOEyv60jmo+185MIv22BfwnMP66+of5N7MOMY5Qsj1ZwKcrgdzAL9FaARObUKstD+WPQ9uE14+X9
eVlzt1tfracpSXRxIJyI62ct1mr4GU/h/CPMEyKUcxEwlrAo8MzMZ/ZnCqPdu/8916AmIkE1fvYp
RbP9jiAoteLmL0iQVkjmm73WO8HOf3EylPJ/MLcvP57FBJcXOaw/w2VT7vgKgsm0J/DkQ1pkcgwQ
IfJOo9yZggLVRAyx3wOnvzeYZgc6sAbYnID943wB5HYNnq6turJmwg64ZwDohoRDnC5wIuB7g1jQ
Yx+H9tSZ5OUYpNfWBLNKqEe3V1LOK5yGccBXQ2Lm01Wjn3QBDH/3LEVvlGF61gUaI9WBsvo5XpUj
tHPi7fX7EgKt0D6jh1/Al/Pl+3UYJhQP+ZCqwiV43AEwYM/VxzXsAzETGHH1ujGgdpwvjQVzWUlN
VvfvxTibVqt8GI6EMxx8kvnJfzDe1ZAMz9y/5Ti1Osmo7wVEGBvvr1p160WP1KqFzNhaqeXQu1pU
fx2iigOsj9utKwAPA5hROT3EpYcGKdTbIN7ldW7aGhMq+9FJmp65vxbUVAoQGmfyZERyHCkjkN8l
UH3aOA5w6ACFvvC01Vm8iEYtGeDWkbJ8wj68yIuW+T+5qMGA3bLR7QPU5vjAapF6gqpzyWApXI9+
IERqU5cZ9txYAon7h9lb6a+2tgpcy5fCrKxZaiBMPUSTu4C4oLMyN2Pir9jHS8lfTr8zNQCDH8Vp
fKpiXJpBj5jANYmqFnEQiVhaaM4KkhCnsWKVUJ9HvemU1oLg/7L6tl6XEN0Km8AIPh9d6p/mVpTd
Ra37ktmmAZnSs9mzccjeSpdMRxvA/6KHMlIBKX/bKKqMTiM/wzr1NntrSP5uJqhxVeOZqzonRkWx
5l+gWZZPQhwKZzGX7gRGimPMs+5NwaXtm/dVqJJZjHF7mVwj3Ip+0pBJHcJ9NhSDBefZmLdk6LLm
kjfOhdMmAfbk+Zoi+s4dQRc86PrAl9V46ypJCmdH2dyD4n86P8BC58xo1S6VVGcLV0esqYuxC0b1
QGSr4abl3OyEnTs1/460xrzpSmtlRIGe8WUtT+mgJd4I8tKCDrucKstvcGk11pY/+ETZJHTLtrSB
14YllpivvOX7UcFh1ubfXhebF9LtOVfksM78QFR/H1TkR+26nN4QIwpTTsSmCieuZtea3v0IJusC
h8H1OkaVotcJQ+5A/NUyFr2CjsxcQyxMbTxUa0OsjiLaD3bh9Tqf9MyL6VA9OFXXe9+6KswN0PF3
s1L+lcQE0a+CXjzvZj0cKJo/jmwaBRNJ4eK/jwM69n8sgK/IzE6vMP8rUrFnH+0lwnFzA/RHXvhj
Nk7IobOdJXnuYHBvXhGx2xn9cQNqQUmgHYCl+SR0boDppVyAvab2MPKaBMU1kSjuE2SPQIz0away
W1ifaSt0hZ9vOE9sRRpPgSi+Hkl8L9TM7X6W3RzaukoT/QBu0hEcmyjxQbEW0G28nHWWelhTbEQf
vdIkj3XBzXcVcXYJ/dEn9VNr18CD4HirGubuJRIBafDmsCqYK28r2nwf8VqXQ7mpQkjjw6lmBSIJ
TZb84188jfud4XoZzjVyuomBhjVYwDPBzk0LZXLl+Y40x2TrbELJk1saetRXbAxVVGozKNKJBS7r
Cri0Jn3tICXzcdGFCe8atQGT0IwPAJQ1AbNyyR1YoQ0cxSuFYPUpBeq71yVCnGM3adX7kpbuMUZ7
gLuFRL/3osa9mFU5Jl4waV28B8biaqUFp1md+9HqFP7Trp09B13nB61rQUsxCrm5Oykk7kh5EpWl
6UK5RN87ytG2x3xhwLF14B3relo1LYs2/QC0Yd9bCqBnB77ein5E4pDmk3LirQC99BaDdLBUeSul
nuRwGQgr2+Hxk/Ek9E/0gC8oxXLsLwc+G3aXQINtx5yZqqoBJ8sFw66wy+dFR5M/hFQuTi+o9Lvu
B/gGcjvXA8DmeZlk7rBgtqd6fr/ax+Hi9FDwtBjcIyYbYqT5i5T/Z9Ct70EjaKQrOoh69abYJ34W
y5eFavtL7WwwtsbK2daaC+cHTdyhFl3UQMqRIJvWbEiKz/WtyBeq3oFNj3hl9W+p7W1MF5dIsJt1
R8eWGVGAjNd3MQZ95ZIzldxskoFd/yoTrr7AFt0htOEGgsaotH4Qdubytgk59JbFn9V7d1Z1io4+
yta2YJbz7kMU+aE1/0CwmauS/dn7cISNgE5/6FM0RZkK7meQRkNAjO3UI3Hp9fdcvoAMlGUdhdNb
l4xkzA3PvDMu9qxh1H8mziYYc1CPH7EKc+9KOJLvHOgptbG6VLPB4CobMq1VwJw38gLP7xE9rPmT
2QtMrp9o4TPeWvY/WQiRD593mZcl91yGvAroO8sH+9q+wuR4SfbIQ1P4lhRVaxlZ+Gw6W9ANY+1v
Sp1Ixg5M6JB5fI4MUFlZPrq7dGJWVH5rGVeMvaI1oYBDOPSB72GHCBprebsw22KPyeTcVQHuZn14
h/PMjmiNnbVvw5L4AQktIjzU1oVpa0Wo/qj9yLabrjBX5xs2uCcxtLAlF5XxuXDLVxRitai+JBgl
/kR1dqic5I0Ml2Lol0YckA5TNyonX46Vr7sMYIbsHX6XEN86n/0KisiFHwx//VWREyloj/ZZYIbE
0AD1EzvNoRWl4Eue45SaGzPFktAV8lfZitxWhtl0VwMu8k77GMXk81kxsYlQm8qgUpZHGT0lypt7
tv+MnhRcYtopFCZrvYzepwMKfpnOOPmQ45ylUcg0yLQ72Xcu1iGJXrJrjn3fkx1ILor74hhsVxU6
6sIZxQcxhTBzsfl2SAHgjz17NPeU6W6Cd8Y0tOP8u4/Uxm8NMIlUw7phBrfu8CRL1PVuVOQal3c4
R+I4l85oCKOxWgMvzozox5p7+bLePUtNChIRj5OoAdmNE4X/8lKLRjdFlDxPr7av+4WTE1GVoO/5
Xtdza5N6CI1KsDQwl9oxHpFesVtvQQviebxgNzgWZqPRtI/A8snl2khdxQOfkvAPApxJzaEAXTPD
QeApIF1blcNFPf1pk4/tvks8jfjCg6a748kHQTC4xXqVMnQuqQ6mO3SrNeSj9e7nLrmiG5a8Xpi/
BcBlZzrC1oC1XcCxt+5qCD25Tv26qci8U+uSSZvXEvvyNgGNZxGK0QEWBGzRGwfOSin5knpZ7rn8
+qdtsvKx0V7CZH9/TgIHi5ozXgvzosUB31KIaN/fG82oUdcTqKh8+X0F/RfYnDi7VaSFaQMYtkuF
rxX9eppE7cOyNHTpgmnGvdTZ73DAW/AeSmHLgGNm9XijnODNEWrMqbBKOlU6vADIpXvzfErqra0b
vGlQnYwBi9sE1MtSRMxB4kiRljkA1CzaukoihCelXal+o6PJOYl2NWObE3hoTJxQOgvm+glYl3fs
jbLm8ah2nvZwVLwdHWQbt+iHY8Ha++7deAmItL7xghUWkYc9rtMmWtsXN2qXAD1hJWe4tbLKAkGY
m1M27SyzKxf6gvQyldX4HMoxYq3YNShT58I40on0uw1khNqfXE5IX9JET0r1zAQkmO9PEbJujdV/
VnrBZeRwuqAbc2/VQZsjv0vTBr6i/t6QkQPppzrwb78dmhWkCjucw19zE6wNruIFXJHid5JMlz0U
GmIFyKDRM9MCq7XUNkbLA2sg24CJWocYkQezTRURaXlN+/HV0V98yeghiLUfcDAlfKl0Z3djs5C1
dvxuIEIBQOOo/AiXfVC4SoKM5lSarQwAX7S+5TrZunt0UNs27vhvQeeHAWnZYSVoBwK/s3FVJQX5
0KjBMXuAzA2jakS8QJiEZHhHxda4uWHy8sKu53kt4vC8/N9QuTCzykuo7pd2WPTxD6ceSctpd1dd
xkaWW9qJMdBTz6AEgZgEkvV4HrVsWQ61cnWZohogRTcWzjLByDFJxML457wZ60hv4nacvj5L34aB
WrAdzz54eaaMicIWXxa5kzbZsPktzJude3og63pi/pbjJx+O8eZc+I72hrlKbNomBVQ8yiCvZm++
EOETBPdw1ECis/8qVKin3bjuYFP6pA9DTO8eY2SCPi3MMHSzwnC3+cBTxuyl3pzn8fYtv3SWc17c
EaVg5V9gFoeEfGP0D2R1Xh50Xoe/eYPn8Buxnxf+SRkidQgZYPtINqI+cvmm2U4dQJJZVcaaEBdS
+vi+r2Jb/kFwqFWovzE4gf9ho8TyAWL8kP+1fC86sJfBV8XxTzNBNNOSpAUdy5JrfjGz2+A3CnZS
iAJijYDPbCTSI9v5jJ3kCjviXDtw+G9IirUJRFd18uFpn9z+9DM0x79Whv1mqzpgvinAbQL6rzNe
O+15JZB2J2Cw7qpaMMvsnEBIIXLAN1lLPyRjrTvqCQ3wbjorOcEWMNoNpfFb71Yo0w/EwyZu2ajo
M56+FdP6tOPopzeRaSUnadH2P3/+ENJwFnQswbDID7bS0uT2zaBegaSbDPSD9xJBQQRiHS05/QV4
nARYkBEynW78XwyQ//srwmr96xRVAIyGJbYm5qIGBL737UOxpg3ib9FXrKtq3dAl/KRpcA8t0BX6
/bbXu3ZIQ0gv6d8/Lwvi2OkVdmkbJ5a/B/XVMxoaG0guAguko5Xr5RDJdNBzty9TRWy42LtJWfFh
pi79WrfEnpB2Xx5mxvirETZ/cVJ/dn7LHy7wJMOunYFR+Qrc+Shg7iH535Dd0b8oVgCJQIWhdiJm
P83HoDGfvClV9TCuFb4cMtIZ3nE9XtHkKTRRVIVMKV7xEY9mM9eZyVUcrBuFDWqyFMIImme6+69q
PXoTL9WGfA2aY55c1cf+vDAF4nRhvxvWJ/70ljFESUFIh3ljhW0NyzHRNXW/uE/Fi9hg/cxV1qOI
UZj311eM1wQlwOou7gJQZAzYgJURmtajzVZIYf1pG2ludXJ9ZkyJqV7GlxuiS1/xJ9GKnZ3KTUhY
fz8TTULigrIOZaXjRynSsa0bFr27OuXHnwYWDsz0U69LcAvqhbF0BXjDAlLNoTg4wuzcfWqoVpRL
jpUVR1AujUJ0Y0KmKJViFRHNghYeCsSW2/c0W/kOEZuhRkUpNGSE5ZKGklvS5QJNBLFCRoz8t8nh
Rmh54aAOgnM2xIJdIP2UK9jbd1f88FZG62BZ0QSpxrtZ7AKr3EAweWnQdEA13MFPrIg8Dp/SBzyb
rKIvW0yA+/BnMuVyKeWo79it1p2SKlPDbdJ35NT/JDkZ8SAdj3Lemu97iSqh0To5lI1WI9jz9d36
Gdw3NSb2P8ng+igJFqkrBt1f+YH4drlmP7dMrMoMCmVU8BylXaxjiiM5GZMltX1vaOVFG4fBbguX
3KpK2HWyRgLPFhNqFqeumZuQrjsXA96N3y+MTxDhFsK2n91vp1zKvXzwJQali7zr8KTpa+F7Evaw
jJ6M7bJm25NhK8lIyra2YMrgPX6QiW6uy7VF2BagrIKGt0ek2YjrJHiwtZOgHUb5HO024sIMVLFM
+3kSgsOrKJlSezOaGr1B6NpygzaAUcd0Vf7ZMe0OOUU1HIuf/C0Bgs0pQm/Jygp1IB5RAjIdt7cT
MVrf2lvJYa2JxRMBbWgv5DpMV0qQWlqysAIiJlE8+XJK4Fj3y1gPFr+xSan6BZf810/HedkSqOFO
5hor9YFFdV96JYwL1kGEv7JxwX8ksZHhnMBH94hr3scq6JoKxTuMLfmC0yvRWnsrPqd1H4mHU+P9
A9CjRTxeV2phz+zvs88Zx9jCBFbHfXhXjOcQ45WcpgiQCvtbeNfeVlUJXg9kyGfh6c0jScHaikr8
zevP48xTC2Z6nzllb9laUoA3fNwTAZSqSwyCZVqXULTMH5V0NFMRlsNiA251BVCx5xmT2jWFy4Ba
lHatFBvbtWtkG9moEgaPELRTjZoZOtTL/GhmWdERp+N5fHhnImzLFJ9lLaqlm+R3DPJF/zxPDVnN
1krIFrRDLRTl/ami6ykwJQ0vM0tA6kDCcxFUBv9EtUeJWJrw2nFfRPPT9CGuxOIb6N/W8RUE07tt
cWJOf/mefk0Uer5yLq+cHmb7bTRNNX8JRseqke0cF6wrZteyH+h4QXLSyfb899QPj8swAZHWMq+6
R/zZogfa1YDRa1pEKQTXqHl32YdDIJztxv6Lww7UcsrmMhnQnzKLdlLZ7QIKpwVOFgXnQlSHt2sd
1QBybR/JA2CRmmT8inz57ujUWZsbrI6uSANBKN+uHeShFpDyjxNE+/gGLwJBJ6stwZencAdMZMYN
ZovnwFwJB8z6cQ7cnqV/HKwjMDj8ppHAiOPJr+vslZqnwiiAhcfzWrU4bgZ4nq9fBnR2Ic/WCY1q
Jp4f8sqtP/x0cj/x3hTMbjl751iZ6YqH9b3S8XxCoHN4T9fq5Z7crMDJcKSew5ekOMAaIPtqEgqo
8w/9BoHxr/IhFDcHkmmLX7JU+knkv2JD1KiAFh7zoHJ+aK0eB3qp++cOVIn4ior+dwTE+qPXf5eC
CAA3MJOLe5tV9ghjByIx50vzyClYALxIEJUBO3rrDGoTOOVHXB63wBqRR968GVjo4l4hrhqg8y/9
aOFeJd9Mu8MNH65ENs6WA1KKG1KbIa6MmudCgaL4WfoOo75tjWvYGM4XvDEjfsLA+StNXXdZUjZG
k8ZvyGsvpVfnCzF+SlnHxrH4eDPj9bHg7dBCe667bfEt3Nh1Q+B9VqRvVLwtL/5OvC7T4nwDdCEx
uQ5oel/uCkx82+QAklJTwfLEgscy+Iq7SsvAHLjojHWelWzG8lq1ZCVmfEsRyGjYgsLUzLIfNDqa
uvYztk8BKPHt9QolZ2Xkz2V0Tqt77nKUQyy0RHmUYYTQSTYksNf5U3zF2c4t6Yl3nIylxgFxDji+
nmyJ9bxjJyxcpnxSxqwt4n2K+tJl3LrO5cPxFqaBlItLEsHfD6xfg++cC1E1bTt/MbmhsxU3VinB
H0j9+ovUV2Lt1rMah+TSMNrEFTfROxKA1b7eGOlChZn61nJd/Hrhf+Fr3TQxZVPDGtER/wtJMR2D
g0QCEuajarHC8B0FcAiVqOEOZIiRfPesgej52yiPl7VXpMrJ/ftZbkMw8T/Vo+WzkaWXFO+USwqb
fkSxVYTmYF6enJ72E4lvH3QwGS+hYw4+qklPfG1GFloiIz+7iB8FGrqUvjuCK3sLpbzoOG75VNjh
PcCVIvJ93m/94n+UyA83IRB6hFqrDmM8TLNX/tRSTY+RLVDInPUdpePLZuNH8YazP8rDGYPhFziv
zgjX28TGc2WjDGxmUMYWBHGFdOJEniAkjZ5XpXCnXy1mB2peI/FXyn1kMNzYO8KpI/Izbpx2WpC8
XnxZKKb3OMrkIyfa9G/qegp/UejDO+1nmXdVmlfNdRtt4CNwY9QaJNaWVJJVmjQbIIdkXWD1YmPl
MEneNIDMMSNYwEd+CqrXRN0yKbgWZVamuzh0NSQ8zM6EIhF80MXHMsp4+IIK28dbWcXHtMEJ0GrT
rJD9eBw3f2rrMNo+0UpHh5y6zQSy3yoRMuUzoEHNU6CckN+S0qm/sYfmWfxQoXVs6t3ahlrcQiom
2wgBBL+ERofBrAaKNDr9Sc1bxdcurnYlApRVuvTwvAAJFASFJu5yYqqzpFLvWYXZXKxHndAto2pO
k46zr8Y00xBKC2DJBuZ5VwZT+YnvduDTdXodnolsWGopOuflM9PjT891AmUgQiLT/1ACZxjTVqou
ABq8/PxJan7Q5gAHJJeooisMh2RQT1lGnaF2ojpsz87UW+ZoFE/q2xLv7Z0io85utf+jM0CpQlcC
GdPp6/2CVv1ML3RPhdadK3Q7g6rabkisr4t4YuEvAc8dNGdSJUsuwFwvXIVWBSNvdxr1oh7LwduS
xdKIygVMVVmRA+rLG6lJs+ml/81GVj2hALymaaCyIjAfiWmb/tejsBC9JASkCMvs2Ecr5hG9XEDT
A2+d1RF6mDju52NojD+HHuq2n9XHKMd1dMnUz53LcynsJW6/hY0XrFN66zPrzmnDRvBC5wtJ1w1P
3f2Zzo0rl6QmhY73vqiAoKQWDE4426geX75tnEaxfevdr/tBKYWsIGJq+hrGxVnlCDrPjFRpxbLo
ziVNi/IEZTOza+agNAC6mBP6L/9Hm+cR/r7vYMr6lgXJAVzsOa0//ktlyfEBuuv6/BrfelKYEXgz
jH9cnOzYixE46eyLymk1AkhPequbbV39oy+ks/T+EdzkJY3cXYuC+vBd4UxO4inY5WmVHwa3qDz/
5j30Ylu5kABa7UTJk6PIYP8z546xo6e7JQwyksPktx0SacS8am/HrTi9gaZb274ZrQunaYsAGsNS
xqWuiRlHHog7bhqd248NFSLP59+StpkOlaXFzt5b7MJUEChEdBiXe1Vpp8dQ4JQ2HB8mQ+2BeXQ2
mWJRRqudY1DaFgnbf8EWNRXyrxrYOXESbrS8IXIHw0K+CVgMtd53vBFCH9Hzo27MoviuJmybKkcu
7JKaeSboYGgsPQQpCHo+bCOYf2tVW+2V1UdzZONOQHZGTqRxtkDYOpMF3z2tsVGTMlhXb8FnjvEh
41JT5vk2sG57/jKVt9JW0h7P6NnEpLnO9GZyNbzsRntsX7HhwKKTJpCyHrqocv7ZoXnz8TnWTBrm
g3x+PyyIKUxHoxthjnpJvJ9gQK3RF4wkErV1F7WHkIvPOZ3jU5LVNMrHOOFnXlMx7jRsocNhFi8U
JdJJAaFTETron/LU8mBEMK8O965EgFw2/3GpFYJzqKUir8gI39Q4K7umGQ0XC1zk6fFs/ngnANKk
xL2bzPrYeHa5jD7YlW3c1nu62Fh7BXObx9IaH+lLxrzFKBBClDmPblrSEW4PnARAB+BY+0AwAgid
XAQPlu2GRSYUaSX1+8AF64HD9cRw34p4sFDIkvD2V4FSqcRjKqGPMjUcLJZzX0LVeVaEJt4/Rzl+
ygGdiVhHsw9zE+kIAOyxOwpJC9sDyvwb31h+FXlowDOrHrLbKERlq0EFnIoNJXyxBAJQPppL/AIn
i9M0Ke6RczjLi6hzmYb/j/yqWBmqNNtsfDa3yGI/wm5xwzBteA9j/qv2oO9E7/jLXqVSwtGzBG1s
0Ev2TVSvwmdWVEU6oPTIeIhjMRYc9V+XxRB6AfkZa91zP7PZG47ANEkM1XVaECSKCGNX8s7hF6pB
/xf5KBIPoqQt1/UzXWyE7kcoUnldMwGA/iTTll8RTA8YCz+Gv2UCbsqMObb5YlfTQqZtzNEV7sLb
cKRkt1gdcdYe2zFlDXROcGcfXh54+xDjIkQunryk7uyitYSYeU88XXjh4lWy+jzcuQkP0rLCatKK
edfKsy3tnbRMXViyo5WpyfC2s8PV5OtWvJ3/eShUnDHi2HaisNnu+qL8FZ2uQBIQkuW/fkBDuenX
i+QXOaqwC2VF3sb/ewWf8QZ9iZwpJKVAlVwjvIhlPck4LYyW2nsHT29AAjUL9Biiv7eT26m6/qlS
lYgNVL5EGKffgaXhbvcjX9B+5f72zxvHyYCrhvValFH0XvMSmisLlwVu+CsQ/VWQldrS4wX7442c
UEbVhsdqO0qB74/EYAB5fUTq7N23umXPe9aPm4XJ6WenO5PzuvFJpBtJMoebb5KUJSr/nAJW6H5e
Py8XyVIRow5CWKRedwakIc02/yM1eo6NVwoODSjEQigiLkKFMv7c0AIgABm7B5Jr9ggpihXmUq3M
EmqxZRuS+l97elsivLyGHOODPT2ZucoLAj2rbnLAwmnDRNl2gcTwVuYLkttiqUKg7IOMqV3m+OtX
wzQFAftv4UpZ3jNx5ydjA4L7UeRNFK5h+Bt/OH17e80NNIkQAW2DfFd4VVzs3yhFuDjWgI/NQvzP
99JogRXNgXhrBlBL3mIDpHrI8Aj71ZJOpjHi/6h7yS6U/ewUktzOT3y3aNaZQK4qrnXfOGdMCoH/
yK8OrYcZ043iVp3QijGQs5VZtQSMnBPwQ2v8lxig6u0xosrl6MqhwKWcZxTah8ee/cGpYRlq+t9o
EU1zDw83ZFcwFXBjt7xta5Ymm7uVWGofrzpHmRgRSx6c6m4D/zpmy7r7UG2jmQ4YMsb5UleF60V+
B7gGAhVK3cWQt1qwTW4nmhzpODR93/CH+X+ELGJbSxjYTBX9htW8xXAM/QF/u56vv/i8K9803h1W
6dPvwhcA9Cfp/ickTjuBRqXwgS+P1yMGuxGqsGgUDNUDpvvc47svXTMXxCIp9ulSVf+NNd5ObWve
6/oCu3JmbQF/VLs6F4J/McyL8hn6hceVNkMog31sH8yKUnXm1Rqa4dokoi5KoQ6a4aHP/beTT97p
PASWuC82awHpMCWmOd1QDKScYDugjUJ0mpoBkVEFRQxMUn9WN7K64YRDajiWKqPkSqVCKyey9nOr
Tjh79HMcj3v0KqzwxfHwRT/WMwcjP9CsiOsD15WaOE2JtutqDMYRm8APgDs4Ypra1D2FM/z3T07S
kZhJgPWqe2PBUrffR2AFrdGZMejox0elw1ux+i4BYaTeG1dyfuGK3H7W7ywYgsyGIB/4KL9K8Bvu
CuG/YEjzkTsSn9bMHbO/1ys8BlGI1GNmP1DoriIYCb4Ldq2kYTMQ6UwzxLxBaa4BwImb6b3rBhbA
PrEV7WyWdXrAy2w1Q+8HLjMyRtsb39tIrz6RQUmNRNqbnmaJXJk9wQo/nekj4ozazMf56aIAPkOv
382P0IrutA77gAoP7x+wFZUyIbKbj0JhsAtJcigY82TgQfysTm2OYkC7vQkcN5Tzb+fc5dElGvEF
LJmewG3Ge5wN1zRPd3JkWIEqPTEoVYzhQInW+t4gRrPm4X54IahviXEAGizHkT9mqCYXcVwpEey5
/a10R+L+qDUpaQszHK62JMWvLtJ3B/XtMX9QHAjcOKRYxDFD0U1q4Ve+8RSJHA5MFlw8o20+O6WU
kaQRYhba6boxveC/ayGD/CMnzw3OSoyYFx1+64Rz2ggLk3RXd1dFidqiXakhU6IqZby5OGi8rO+9
T1YF/mSHpm3tZFa0V+HDxeblLgbC+XmOWC5zQyX48CuwQPZSQgYaTCqfdwK1WH7YkJDH9IHwtgWv
YXj1iVFhNNveAco3D/VcCjUX6jpaA/pAhLyTAcyAnyYZzKsXFSjH7Cf60XlgEfudK/LRwdXkE3ex
BGF/95ICbrEqx1n9JDaaUqitb+2W7HtBCkhsAXklZYbbeOm8Tiiu9Jj6goVIFaYPUGNGf+at3ZYJ
UjM655Qcu1FOeanmeebSi7zHv/jTx3lNAWi04pqbghRIgC3Mb8ZZ5saGWfePLL9L9bsrYrLTZCEi
/k0t+uH0QbDMKtm6ihat1YR/NmT2hflW45GkNqIxyHgjLmncAvhsWNxUGmKyZ6Xs8phznftV66rd
ossuF2+Q+5hFtT6t0iotaZsvxxE/HA8Yv91eGZJOM+UtGk//hvOuBIOA8Bjj44lccagW7uEDa1Kf
3STjVZlKjHFF1YmUp4XW/6Tj8vcUY2Th4KacCRXAiByKhmO0Xn83oZCMfCgMTtsEi8RgQLW1CA1u
3lcVKk9Yp6L/xrsTMWJ+PdRQu32uW4EgA1FocgxFbN8Vj4pOFsfJ6otWPTuLjGyexFDXiz5DNUnn
1DB5F6Tmo/BW2oEVw9jdDxocLmOUSe/PXt5Fzd2LxMhdVDd2F3JZoGhIZ+uFy2hVQ5w8qSdjFsSU
4hNthx7ukH5pMBpp6OxnEg9+Vc7pjK8dwwyOsk2WKDvVECi1ovcDVGJB/ONPz0BWGrziMKLKjX39
tjnugT8w5Hv+qjT7UQWhlkynBppUvMtzTi/l8RhrVhpwbf+cYUIRjI4mbp+gv109QkZN2f1jEd9U
bvIaJMWggurWpFwVezzBKBbXOJS47KD84xTp4q09FjUDzAtbJyiasRvteq1huto029EEMg63HTPH
Rr/PRk0cnjIZHvZsUF6gpz9J8yL/mP7pkq4dG3J0KzxgGFvWuo3B1Xb2+CI1zKD4EgsYLV9z0yxB
wzgXh9V4P0cBPFOOFvC2OAAlS+FU5xIVcFMXj3Bcv+/k0qt3vv4A8COIN0mOA0LYvu6/jHDsmg2L
QCXNxU56wm7bWEGv8hr7ZrE3GKX8YXcYWtNj+lKHHch3EiE6mZpZvUzyKVAWV+kCm484HQe6g6Ba
GWGSe1WNXXlqn9Lr/e/KpzU+LSqzjUYNqBBCPaBQqpiI+TLQChoYeIdUgqVuHthWJ8ZBUGBVYvz+
rySAoYvhdgFQur4rmB5qv/iLlGV0RsEznZhrVpJ59ey9iHpz6wZO2bxzAYnO3CUXlKqigqLdSvOS
wTm/bdWepciJjoEG7L/4h1iTlxTHG9ic/Z5tCspJ08KSxBANYBCtSXtdmiebNfmFroXw/ApLFGEo
2Iynd0vL+ofzZjVAHnZjRfOtnkY7Knzb5muukIrbNRBcDRgKT7/Gn+k0blxbjyjXFFTdJ0SjrXxH
V6kGhqgzibVvHN0t48CgZLEecbI9wc1ZlJ/W1pu2eZCHbpzZ6YS8ubehig6C7KCa7r2TCS6NS/Ua
O0gEK3h8LAV5qAmTxwqqYUZ6uWWiD1swJsTjuEVhl6M5iog5QeZSeKP4tPt+1Kt+qth3P7aIJ6Xs
9hrvsxRWBlLjfKfItsd2fyFDVteJ5+hyXfWGzROlVpnjARGxp4KV0UkDYRpKjo+zazT4Xiv0VAnp
vDA25+53R5d/g0V0eIFKx5Sn6K7GdPAJrmS4WD/Y/iD6Yfb24Pm0pgqFx8NwFQ12x0ZRDUy/f8To
Sg6QXHpUAEfGiPXIL8aLB2F7P5uxd2MG/Pciu10jKngVB5BKtX3L8GdRJqhQTD1B14petVbwTs0c
oVmEWgnk7D0565RspyS1+ZLfiz9ZNvGlDpGcqOj1zY5XFMaGdGv/rQVJ+M58MUrG83H2xPKhMfHB
U7yGHYpcBnsTnXkNtTtJablBVyW4pj2QlRkycjZwshfk4m3N9+rT1C2yDm5+mhWxUrgY/B7OC7KQ
3+OwKOvlhj+vS6IngWrIbE8CUKoNQw11pDYmFFSA1M7G05IGchhcVRJq0K/ll85SpU5ADDqL0m0m
NLAtp5gtWfRoOmKmlDmZS1h+eGicfbQykgebEl/jeuchA5SiJJK4cwb3EKqsObB3JSK73otZ1OIy
WFwQgUfNGNlBGrGVTJrPbjzfeY8z0UQ7nBzwX+TtxtXpH+HRlE0sgGS44F8OqRcZkVaX6hqoJFJv
Zm/Odtk727gPafSKAYNwQKarNMVdDbzN7KH1zhbUoo5Iyj8Eaq3qpge6IluWuZOxN8hJePWOgnwC
nogNWrMOneY16THPRJ+E+ucH6YchtvYfXeQUeaksrLcwRaIr1If9/9IvxTz24ZgONmfRh8CXWN3i
pNbGmUSas2th9Q9kTF6gKtCBOUoZOB1qGip+/TyXTvKYHj/BPiHgUf4HTyLfHEUXEcoWUYZbTcqX
2n/IrNwcWSUopaBY23w/oB3qW7mr3mUID283H98UPEx1uD0AUnwbx2mW/xx3Yvo/kne3Cv3Ps6qj
V3iEw62pVbZic+YjaxIxp/UTbZ2tYIztZRV2RjndpJW6JDouTir8iUTH09Q0HPGW/ILjD0/AKdx8
RJNiUtm9wy92aniPop3IXYKdTpFhXy+qPMbLT5SBhW9M40+rs02X+ixqrKrDk7PUqZNIRS/53yKB
R8G86UluVkAoKM16tF4JulluF2U3/TyibQvadrU4y8B/noFzMbtfCuJonSb4xb9eANvsry91IHxo
WfiL0E3t7ehdo1/6dYeQ+FeWhd1sm6M7sZHjfrjV8anFIjgooiDsQUv/e8aEbqAt7QYg3gZIJu1r
nYsANspL7SYWS9l8YpcX0khi0P0u7cWlrZQhGVMW9L/VeCkB50nvZyw+sOfRKRc3QlQ2vM3CH5hj
v0KhMRErqOABK3ma2XvZN8cVOqokeK1ZNfNK8Xjdt4IT9B29Xgr5xtNnJFi62k65Kp+DZb5aMZtd
SOLVzoi31QU5KZBDQ6CpzTlixvQ4lIsZyyMNXSDGyW6IhwE78Msm8D5IlI7zGOc+oq/ZjfD4CRcN
mcQgiltXKfTwsQmXkiawIbuuL6ZKI936M1iw7SXXwJ+XybpK4otjvvJdriwKRUBMFf2bt3rGlIrD
VgWfJNrykyXffAbC0DP0e6Gk+ZdJTCKN3eGJ7N/kNNW5YfzKneGfgkyXnz1ZaxJCv5OJiqTma431
VT6k7ec7UUSBX7OsMqhwasRIMn9kDS8d+b227Q/OPxtQ3hntvsJWbZ9ZD2DNM7eOXK+tGkrbDN18
Z7D9YtfIVYX2wcEa9w7S99O7OEcwl4lGt5dr934F8Bf6g7LVv4e9ppGFpq3Sdt3tJnhp/VyeMaag
zYUvZXHfOSx35U3CujPpLPU3QEmDgsgY5W1fpOX2zJDOYmto/yI7x+RPJ6mGrUtjQSrbzuVQElHt
ZzINdSMXIiyy6iCldZm4U6QX6gcRUYlpStmKQC/qJv4AdFp7gPR/ArX6x/1mPFn5J4IFsJb4bfZu
hkoq+UqpjkxLQ4dW/rEvpMQlkKjnaVycryapxLVoKE7xUzRP9CT96BwRnHdSbYcuRPfFotpemj7p
dAUsqNgunf0SGXf2N39UB33KDzoR8jRAM1UVo3TNuUdyGxQjf5X9s7zad9ZDOXW4fFFRLeuk59As
XsX6sXIb6CmJlzPr7RF7DqK5v/kDXdLCEuh+xFYLk44fQuumR3buDbJXcnqglULNEyLBUCw3A9r9
ZlTnqXuDA+EQ0jPXYEelYFGHp7gv29LCGH4GOyXfpkvxyYfcVJgyaz5wlu25JT9ry9WHojOJBvcE
c4CDzloXXrxEGrE/epxyc1sL3XhAtxOhUYuK1nTZultaI+ZoQZOXFjhEOrYzNQoKnaUfyXBmvlzS
wyAk4Loot6ypNbW1LsUtSh91hCTSLs13o/kiek/RikqoMo6HLk+j9eJyFPAVoyH9EAhVF8TEFZUP
YYwJqV8hjcx28FqExo5U7qq+iABcqx3eCjP9ll5UTnL6JjMDCCmwpbhTU7ImqeeDFIW4WJPr9VaX
5iRadsF5QrkTrMiX0qdL/QB4OyvlArE850/uZe1N+ktXzhJTE9OGIzaQzCqPbp0FhObwEjJJES0/
pCBb5OmP58I1k/asstcgS+oMjNo68ecisK/3u95ik9uwcRuH31Wge7KUfKwraXhvcsoGniyZAq9w
cRqSWNWSMrPh0tcR8A2ukePbh9Q7aWBGABPV3ZNmvdmX0e618+/JBKk3ie80ERpntdvAh4Qtc229
Usem3NLQSQCnMFHBlfuqKgR05JHiLdymmXEAIrRBp+PY7a0bmC6bTN5q7LTcQZIKEQH3mZqzw11O
oopMDYK/Rzc7NM1b5HIwKD2Qp60X5TThXgi5nNXTccxAWgLC4my6Pg/Jq+igTSG+nfm8R46Be7m3
EW5Bk1FBWJM4GjrYOxILH2FODhTu3BL+QxTqNWTYlQmMBfTNYhoG8pRCb+zHKS5YEjRPZs99gfRe
crADkco35qinuEvkd5LwhjqkwywafipM0hJGe3U/C03e9xMGWHSNdW3KUqADYMo+nuhgGNp7VX4M
fIUrvBsBGyK4Brg63tZIUhUat82cFmkTBQbkuV6KNjMwS+piX3KAq4pqmOrwG0JyJz9kG9UKGhGb
ayLnsIf59xDG4ccHc3df35cCLQNmwzSYyei9AZb6lZW0MI+cy/Tj3Qv7duMyBuhM+Ef/8LwGuJ8S
lvgm5mlkeo9bZyPD8TXTYBKEDz2PxJzXBdC0c27tKoUnM5ID4zcTN0OnUSHQ9kD+zz+j50Z5y3sV
5OHyjmGd+X9J/BAr/+2RnoEJzi2UsBh0ARCl+hJF4L2Fu13rr3m/tmMVElFtzmsb2QT/Xl+mShWS
KTUC25tA9tIwTTvn5mKiXQSWIbdwa98+S9jE0+XcnEz0S8aKpWPtDSZbA3ScD3Si10Vu1WhXNbEd
m4viPjuYaWeuk2xmKmvxygn99jfMQLibZKVZ2z8Ze7Z/sQjrElBehdQEKKiZ8RZy5in1fKOfA2f0
e1hImX7suGnKNJuGII2d/HyGZGCs4KZFVSW+d6BNa0Dmhs+LNtZN6+3uVaBpx1GPZvGReaHa08Yp
zucorE+rN2FGBrdqLUOEnw5BszkZZF0m58W/sUzIrciyLWjzIcZAUYRupwL2VRhrpIV9SA+63CDn
pHpbzm0/lOEgHRd2ufuLbO93U/zesuJpbyNHtAAt4ZF5XxogFXz9LswEm+n8IoZaTzqAEOsSHyu2
kx/7CF1SrIPU/lWPwWB89QV3FBGQ3xiX5Gti/EsDPOg6TZiOhACiwumZsnWixMajl5sv+zyHJ38h
iuyRxOf6QxJ2uFLPsuaBoqmB6w7RB8Gev1vk4tdrg8SRSAJlMGtZGD2vvipKzcvj1EYmGqKpOgUB
oLMaC09Wa8+Hj20SiPF5atH6Ddwiqx9HQDJUJrOCX3Ox2hcxvLno5WDvID6+LmiXLIRLchVIzFBZ
h6IPv3WkQ5FFsTB7Id9eqs40N9PrP+bH3nlv+jHzm+VhS+IiIw1ffxmu5q+envirBuQLYASIW1hs
qVtjjwr3SBHU4qTSR3kawYjnVM9rKfiUkijVur11TeMPdx+GNWskMqpeZBP0XvsaWPb0wGkSnfK1
cyyhGnTG+dfBB+lgt/vXsRwj+CO3BBzUVGo22p+vCvgRluNiAd2CuMHbhe0kjsL4RKgfO/SjVo74
mkrp2Pf6W2rlcoKu9Iu0MliaueNpFZSHChcCehMsEyznI8Zgm3TCpdunJCIt7cODbExy7GbR3tfq
UR1AwK/RpJZb0ts/soneCl/wpWfk4Hs7FgkNl+scHIqCv96IEnpmbn0JxD4PkWBEaAKhMb+jyakh
kKg4z6lJ0+SVLnAk0f3vGUrNcsE8wCkP4i8Ps7w/he5WYrt+DIZo+qv/Ai/tx+IkCnVmkzihQAmK
8rGWGQE9Mu9Gz1utM1on0M1xDYGx8zRt6Eym8Dni/T/mDDDkyAPJKbPngFouuNswtu4h6j21DVnB
+7ZAZweICGZtWLhNPvCwH37wfnYoYsj+p4rmfRM3Vml7EBwoB2xoPTHjyyo8YSQ1YXaTXyfElvoA
fRc0XEnaqUAX0rpHDZVaDuB9pcbBZ/9xYpLovnliCWKBBbd+7mFnIW/LCc98TlrVydJsJWCfZ3lo
ojDYwCAuzEQIKGZhMK85k3M3v6X2SQAUo5ID/l46MoEqcMSvXpPQ6Z2ZVt9B/MrAakg1jZM43+bC
5YNgsJMDZuQzkZ7Tmh6t42MVW8ooE5T2+F7mkIBsYWh3O57CjxpVhTSMeq86AmCDdRjatp0sh5cL
ptZ9+8fGVG+L4wyPWNrUlfDwz6dFlJsJG9ENcbnnFd9QM0uYN8TcLZScGLaFVJmSXdy0UfgJUoXo
MvViYddSHv4Wj9jZyYF0ephGJwUSvhQTPqiXAb5Q8SzIGkfvUtsj6UycNBJBSegfnXvWWoZCJyeK
ZTu/CHsOAu2zFR31Rt7ZDvGyksifb2K0Q4Lk5PMafunzciDjT4A7pPjyyBaLb4mbS2hcu6q6PkUT
y4HdXPIzN+yYGEslRm0OGPgd3chEc6X9XymftsUsO1I+qJiS6HcNCx3REazgyrNTltZPV4XfRzG7
8pZj5EnmoqOiwRU5S3P7rIFB3VSec/k7h+imtcjDWnDwnCEkLFTUibGtFUieRMeHgLGrkuW7MuJL
9Zod/TLbXiqZe2qC3ZqOcgQKh3xKeKoPrPyObxcLAr3zjLscaac14XZ6mJO71R/6xWV23TUbNLCG
zFVZ2HRaQdfC9K+kxTf23LXRB4cCtdmEbc/sFTHQSJKukUg/+QHhpUsn2CSrhUam1FHx2gomRYQs
uUcPP3cU/QHOTGgYFyJSh8FqEtYOHDVc0XkFDH675NDOkbxLXJ+tNWvoySd0CTfQKzj6w1ONjZGt
SoWZ7hMuP3dT55G0BBWZhw6yQA+8gyC3jqPmjMmJ8NR178+2A23svLKJ0dJXjR2voNckxtOFVB+2
G6a+nxndSYJODL5HxD2WW4iVsTeLPUTA2It3AOIeLEkOA5p5i9/XRhaqRgzkaPSfyZVCutI0xxik
oqVS9hoHtaIHg1zcfzt68fNFxcuGc+MlFMABaDq6uiMqkrLpOXm10S/Q3GUwD7Jqb5dKVeu0bmLO
nygJYIhvEEG8i1Gxhsiop2Fb7AouOyj413iOyqkdXayw4WlSgHichfAq+JEAr0gOp1n+M/g84NtC
BZSo8ecVefUcjXNjEzq3/nhRplYiAR35sQpI3mSFiIaZL9093m46On9I7tDPYlgxxkVmA2zdUpJm
LN/QrFI8Nhvuox1rTFf1ZWXMEkS7jr2Hx7XghHPRdcWl8tX+u1DFObApFItl5JGZeWT4s/4kxrV9
MZYRKDVeHsuDPAik/KBHDcLk2yk2jy0ZV7zfCrVvgL5lJS35fCfeg6Lf5hvCDevP1/hjaL6y6GWQ
aI/qs05vZCq/kFvoQRahyW7cbmbUJsi3W0rgX1sR7c6nXEPDjFezCUPXpQSLi5rObwT64n8gEV/5
MUNGm55y9QUVSrQ3xeAzaMSdx6nE2QznMJZeqMorz4FonPXCJPqn7mqffvvnmWrCviIm5W2A1Nnl
PU3wQe6TZcmP0CijZLUBpCVwNWhzjje+XbncZstqL8D9oHecv8dvbbxKa4WzcgJYtEVLGI9Fm9xs
ytsNpbYbHt8dHAJhRzuflp+w5JJYq9rhMu77/dEPuQKpyXlEL1+YzgLAca0uKkTkp7yV+LZ85Qbg
r7cz0MuyNWhYjsfZ1A9US28tMmcUgkHjs+pZgNjNkwJEVY4l6r1VB717Ry4RWblPvXdkqHGfugHb
jaKtiawEUA4twRjLi/bi/I+OlfJmgrBnwCQRxyFhcfr56wOZSGFTuA7f0i4YOVQfOEfFuKleQDP3
EDL/1vM/C533+F4znsNbGP6oFLRPyEloTwQsezR5yHYBhy6aYRdG455nAcJVsQuPrhORWVcmloyA
BtGSrg8TKYOg8BOdd2UNKEFmfjicf0yLbpzUCsK+n1M1d4TFNPuyu6qoM1D1FkDCefzckB4WhQWz
Wv2CLAN/CJntGpykyVKx4G2VsJZgB56uBIgi9UyXrc00ByivkIINw5CQ37/wwCAgvdlKu0+MLRb8
LdJcm5nwsAk62xgTQ8TAR24piTdTZCNvI8VTbz+b4HcR7vuvoQRvsmvUtkguDNMQS3ofIczb71mM
EoVOeJ92Utu4YAzn3mDEYAbITKAJ6prUgn6eBIEOJ66+kw9/8SVUVUl7rPRV3vJvkizBOF0Acxq7
atBcqDteb50l4S82X3oHxe+BNObQv9X1gUk0nM5aPaqqD9m2OMZd+WxjRvFJetn6awk6qNk40I6a
H3Y4ZW3c3VIk9Bo4VAtCz0U2ZfzkW0bdO87cvoryvw/znsf1/6Dqs0Py61n79YRvL23SUUQ5sGaH
CWK7Ks2KX0Psw+CjYdvJkiSIqO5A+hahk59Oztc7gjb5dp1yknyON674MnX7jsTvNBj3qBCsg8va
aFB7MYeca9SQ8a6hDYc/isNbFDx+9TQq7LchUpHrhvhwBkAIfhQ/9YTolrd47P/2t6eM2vlV7JCD
iUIEd9cz3yIe0xOCs/tf6FNYQjRC7UMwLIKjPCFPZkEzTUM9QRYJVgNc+5F/T+itLxmkk4jpma0H
BzqRlI8ErdzR4SQkUfAIlimbbQmVx+FKFuOYtAberWMikIUFPMft6nJ/1LuQj7RlYknfPfiZYaMO
bKYcTfrSZgpz+/HhNXaYeOr+w0bTa3YRpFX1SdxjqoiQNQAqv+MTU4g+yr7P7esccVI2ujzRbHKk
v46HsOr8G+6KAH8u7CobRnO/KAWtsce9MNk1rsEDeaCf2b1nGQiaPh6vm+bRHyqqLlNDf2zHiT/R
iLnI+/29LUokgi318LS3GC2yuDNuHLJ8b/5JEcppMrSHakmL5BZu5q7au60JcJeuf4sFqcsF2JFS
KrtZjGQTKd0/eOHJjF1tTW6ZCcBhDHAW+piU9dBrUuizXRhhsz4grF0FVZjSwwe4Uw3hcUKZZQ9l
Fzv2WK3ZKUa8r3PsXsGyRypb+vJ4/ib8S47w3jI69p6U7cVqgWSfb5AHQpHYzfxy4j7HiQC2rFZU
1OrPAC1xgk0max1UfJq8Of8ImiwDlV/CEmcPMHg66Oki1FttdFc9hPOiQdH9CSuGBLFbf6tmKFl6
6pue4UeKHCV4N3jN5dlQMs7EpvnS2kSvj7yxeMO/vv2HeCBoWXkv5uZ2KWRNEla5S++XHNkdDeyv
5PPe1He1OPVlAOM+3vkkKzrTlZDvfb7lSr8257a7toM4iADbUuU4rMkuaTK/XZD0Xa12TATCrLrW
BYf8WVeYwNnZXaDsJ8eCxTZIZmJyBXSKvtx3yIeOoc4/wKaWfAzadR2xw7ODU9O6l70GEUniiWW1
ZKQlZjcSnvNc5putxDul8uQjV9I5O4ZU/Q6CYLr2KMxE3adw4fzlTRTpktbOPZQ9qSISajXdYNEi
vKRVHAgT3qD0Tb/VUeughVYgyoNqL9q7LINArJMpPIHzC9b4KEA8XROSlVFQPRacwDnih8eAbyor
FHDFlgCH3ChRTeFTxAxsolhNTERMXq2kA7aqJByyp91oCBsHotTpODlD70mxy1l2lCRwKYwOkO38
i++hhSznz+IofylZY17qfRC8AxhY3MJyrSHbH9Lj/yD40ZCKUg0SI6WmU9S6lgCADDF/8U0iLY1q
UzxhmsY0oUa98z7CeZiiTJ7W23H9vkLs3uvK2iVJ0Zati9L9cViGOhhVbrjwpB03n0MEUhRSaMN0
YuiXnpcyKnoe9Rwy+6eki+E39Y0DVh/wRT9203b33EjANaIGcc0ECJtUXQyMMTTgr3sBwLk8/Ej2
EIp75DksQXpF5ASnksYebb18AaQDRSsRvcqDQpipZcpbIjsai/g5dfPSWBfjFGDPvd4GX0GxFbXB
Id7YOl9Gcosuw/gsYRpUzdgjlIfJAmpeMpc7mUoH0fmohcgSAD5X+mwUxrRMa6Lvja9GZqMgQcso
9YidstGLgQ1ELlIy7cQvJwKOCZ6Zapr1jAcg7hD9Z1RWvANHP+W35xmKz5sklqRXb/rp7VV0f9to
PfBo6g6BP81fMeisvFNaI4F/17qJAdvwTR0wPIxJkRYGQhjdTjF+9HP96Tpd0TAlwPW4qC9/ySl+
ALaAKzKK66/8WR064MIIwSvDS4DcGFfAnAnbD9zfbeT93P1ULv5ZJ22roYb66Ki9ZpmErZkm8FpJ
2qyzxL1M+Nt0QkyDXFIcapDB9HV4PCsgtdgPnwMfSbu/h9VZkVXUifHxgQQIXv03fZ7OYQHgqOwx
2RH2wkle89OEncvS3f7RwW8tU8gppIwptvPNpZrSbxgiFN9Pf/be6tgXshyfNi6ywRnYID66WVhX
h0nGWx2lKFWUehJKLhIRMG538THGZMif+b8NEaIlrj7sMdUu8S63oJZNgWecokASkGcCJ13VXkP+
8XML/39pFZklQcvgjY2cvwXZSrxrQJfbP+LFXKgHPeUbtAxDCHCl7lyQmaaOMxVH1sw03ACfGENf
963mpLCMviGJleJvlS3mylwJHNZ3ebZATiNtdbL3PQfq9y6WmAoQPk161SCSpVvNeB53D40lOF1C
WwgXlm98+jL8ehH3XeUVZrLaEEj/jpBn4semZ5k7SXHe6PDK60AW2R6hGwcoXzimX1E0uD58ZWcb
2oxTgEXiyZVEy6iwy9gM5JWqKj3xZ12xprS5wAN7Sdu3Snr5/kgNvB82sIk97LJ6+RZp332POteO
2fj8P+aqnKHF3WtPiZJx2e7S7xXRQtE/ccmE51VBAT/kPB9AQeZgpNufqwHFYcpnTvbIEtSafPEz
EqLjauFUpESOlV0eUsGc786/tbbv47n8SmW/g/xgvl6opTu+7jjbKmdVHVCMT2Xs45NieOjK12aD
n3OSoS+KIogPDkC6uA090TU8TcoyO/I2zsk57wRtywQgbqQZ76OgO7uK3+msCS+vVwYWztpxOj0e
4312QuAdfhOezvGhOJGwMD4w5PumnAlvX7JKJ8gJIh8Tp2QlGhuZzMns5SV7DTcUEuSJSBpBzUGp
G+s4nt657hpCZhOEYsa9SdmL4y2911BGE8+NDM4sGun1L7qYCLr2sc1WDTAHN4UVf1TqCwZ/iNGW
+WxwC8oE3LXpwDJox1L6KxEVZXy37tzRGpF5ER1CNOeWoUgnNaGlBaJdsYXoZpMaguTxXFEQ2h1A
FySUbczBeFXtvOIfyYohAjPRsV69NP1EpWf1Qitj1q0Vv52Ka0/zpFvUkhUAco+3Ek+XzZAOQGYV
TpZRmqbOe/m3HndVR0sFu1D56pE3ppq9VDC5VaXMIX+ApD5c9GVVxAFm6agKAq+/Iu9JpoSJ0nr5
5F0k9QQ0MD6QGdDd3QlfZE+BWRQmccLyN6Ykpuh5IRk86MMEvlQ9j0wRHgOxusj2jmJfef+rD3ph
uyb7NCSjIX0NvuO1VHnG1mkzebbMH+AYuGMJZ8PBmkG5x6nIE/rdE3J/6/Uk9m6FTfM6jY0TtDUj
45OUddGS5azMalR9FA8RCuyg56VwNMEBCcNg2ZABCJfUs7aZH+BuzwlBAMV1GjXqmFGLs07KZ2Sw
aFSFqzecjxFk/HXCwYUNS7NAHCSwRVgsPeOrp3yZOOKY1Yo7IjxHG2MA6+0m6S3p6WWMILNZmsEK
gXTZswmN+qDy6wUVXVjQVQ6ZlacVRg9lkt6ta+cBNcHFFUoftl7QldOhrYLwJPpgRvHdtJURimID
rPN3PdgCYC5nggU1POoEEfqxhm7Q21iF5vARZdakc3cVSYQa9/Q4FLHCE6PqHipXETxeZqHiONkC
uetpbhki68oqTMiqIEn002wOAS5Ldk/Evk8yi9IK8PdioLDGdyL5H8+/wvQ65ekTeh79/feq3CsO
ivduCAhZytgt3D0szMb5k7GDL1FzgzNUrXV0SFYkryKsnklOxeAxnSVAei7pxdfVkwsmsSAYSn09
USs0RppqHplxn3VPTVwM/U0N+nHqsrb5uy0MQvoxyt/d7U52xdcnub0dJBvjodwOYss9mfP1VVCq
czBrS639DooNjZXzmZOI1iyiZzIyc0rx+kqBBm9xlVJ5fjMmKl05KIsMBHAwR+epPUfloRn+Z67C
w9JmdixTiC+pzQPboBvKXkcZqnmV+lLrwbUIfd5Ejdmdw7xRAdQstwes6xva11F9oI2lkgrlQRHV
L9FrbRomGWtzG0yU4Q5H9Zj9MdspZ6CbcgIOEgfXnCwmmjvpx5ftdQldS4TjzNk4yC8jV4MlpfQ+
GT1bm8839bnrOayrdaDy+yS9xUUwmlR8sWrlRTE3QntKpD0H9jYPMtG2QNlAbbtVD3tgog+bFiSX
QWPJtviqGUqavQjxIPRU0ro10ohTIHyv8B19G0iG8I64Ya2vwT7mQqiAToTeMjbgJwFYteJAH2Rh
LYuSLGQl5SixH68tuedLTUCByIPvAAtwWBX++sx5rJ4HQvYcZO1aQvtKbKg9Ox1IocpD2Uq0qbDs
3VzkwBqO/uLFuMPprsWE1MAq22lnhz15A2C1whokhew8hStGg5XP+ay6U2VdoC2kjpWeZvSci0MO
JExO105s7PVLC4v9H+z/i5//ck1FiZZg2hwwoB3kjiZ8wYx4ocOeRBZjlRlrayS0t/6Twehcy4+J
LgXdY6dgSTsY5xq8Dca+p+e8VRPDF93A5gCkYsZkQkUF74cwAiyqhZsCip3mLabCtEXxEga2x9+W
9V4aIVo7z5mmVmE6JFyM/DBsWzFfQPX1izhpiO1S/aywTA+lr4Q/qqLGKWZz1b/fyLtVb45ko9Ui
q0zt/Tog9Z47IbPjrzq3fOuZCOa/65evCvj+SRN/mFRUrEf4zgipE3cRK2vCB47jK5q+TZ/74aay
8epWI4FnQgqi6/2rj152GyAWVMDBOlf9GpC24+A++BqsJoL1xEul1SMp4T/JIs5/obj5XBMocwgr
fK6clDGDFFt3SjncL74XOoxPHNvlPD1v9XnrV2/qOotVgxqm4gw1iuLTEQGDtSIkYkp4NBYdJIrc
OzWFvAzwbv26iItQ1WUcqv8bhbkzD/5IzFo3a04QOtlwydSAbaEx1V38oOce+3npHRHkvV5B6dTU
rzhUSfg0bmElVH/C91Dnk0Qh4njqJF1TLC9j0rknaESQf8cNwzFUMxQza5arcgo8HoWAMZpUUGFY
y9d7roRHmX/6dBc0j7UFJDq53EKSTFsfXjBRXFN5Re7xUYTok3VTIzrQnx82fpfxiOfoKfEK0r8w
qIKoifLp9JJQcK5mXseLtNkVWWB7PnkKPnW9ufuRWytGA5E/XEVaAe8giZOL1WoiwtMof2MR5SvF
w8YGtirLqndwb1YhHKPQ9VLhW8cp5h25Vf8hAqLtgNXLxbrUFH7Ni+pmnlof21Qai+ScG8H/yE6F
3oY0c9sCMLjQpIQhWIj8rPzh/+FVhI21SWcl7RU1UIIQNaJOQwsH+nbhWP3aEbNpaiq256LXgX4Z
syhxfjDR43tGHsLDAXsJTG0szPK/w2LDMJaOkdON61dpEykUgkCi/yH4A1GZimtpvpvKWne2cnUE
L1/xiKcmfFi9745DlZo6X/ekLMA0ul8QcnTxTtMRzI1FeWi8ebzqfn4UZdhRa1E0o48LaJP209GI
N9QCyi3028Jb/21VzRy028sZ4nBw4qID6r0WKuep9dY61hoteq6qbSzicYmC06lHo3wfc3y/vXp4
ts/7hlFRh+sPswpQ6LLS01gOauf8xE6AnUP3Z03PUJuSRleWv59vbu2vNSHAzicl0FmWMNQdFQKG
x14lHE4BwAgUZVLisw2xhEV/DmTWsxsONPSJhtcojkfL4m5EsytMcyyEFfSyUL6RnIWQlIxcE/cf
o8EpshMWxBuSomz1brEx4ckZxN8Bsm6ev+PV5wStrZOa5kIne7DXt1bI99ri0QpfdzSVoFdHObP9
bjdAgA9Z2GeC+2x8CBQyhLhM9+L8m09pY4A2NZ1BX8/aRmToHPEN5IuKqjBavPpgzLRozeakZ+aD
/KqZ4kxUxdgAmPgoEH1QZCkcW+SVJJ4PRTNIBra4sYQwjbzamT/9kq/NLsgTZOpIHzWa/WrWC4Vc
eKBFBlWFb2CacsR7uEKxCVOOOHNNzKmhPUvkz3l8Q9atX5rd8Jyh3DQG6yY3b1bh8b98H8qVxTtT
yyScaDUCaxz9ueaKF9XM06IsNB+lu8uycys0ZdPWbSCDXYaukli0T+0iwSpJIdUybSr7Canf4kyd
WaxK9g7An7F6Mt9fBwUaQ8dSk4yYIzCyq2TTJZuJQhf/Ju+lRnyzpKEefy8zt288zItlebUh0EAj
gercO2cEe4yEoc8rTktQIsa7MAkBn4JYILr5VLF6Ksj32QSJPRsQoKI7NqpcuH9bJAYfkwlGe5ko
DIaecJEXDF283hmi5lNOAFRe6QgvzNyFOGALBGUpIqONRGn9ddlkVcwP34b1FHoEb2oel7zZH/r+
ocxQUe3vgIfWx8zYBeutkGOp4au2wrRX/DVuwzVAZ2Z2C1yfxN9utlOb/28TFmTCuO6mfZM0gezj
X50DjlJ2fLUKs2xQXoE42KhRk14KDjMP60bCfWPsr2+gX4QwhRqybxo2diP7ImK7+d/NK9YFmU8C
vXkhLfd3lNJSTSVNRlLluuOj0cuMk6QcrePWNVeLnBxpdvIhOpbVjU7s5x4+cNf08VZWDdEyZPuA
kdNKfCC8+6+0D4BLOQB5H/cSBT93HkA2wg/L+lj+sSlCQGeTAxi9dKAOZ7FMpbgI7UiZZyNhB+tD
vLHlWFGzpJ5059Qt8ntCa1bhpKyQPudpajn4bCd1gRPsm447oWv2KE618HVNYXINEKv+ATjHpnWm
0zoP61so+6wGlKXpDFvZnxmfGlxsE6z0aQmneJ+Vr0MoJd1HhIQmZo5wBjcSBbGzpaITpFTy14WX
c4w95i3rFcFzOVbzTq+57EFTFoyvEeJPMlcuf/wanL+L2G59Y+5P/oih7mtSFwbFEjqT29STET5Q
mVm9lMFbjYQhusgDdh66klfmgmc/cLPQ6tslsdTpqLyoYkOz4n4IJtFBoVO4kjn+hqSzqLtZYynz
tnaMBLYYxr2gPu/G1Xz6UBmZtpx1emp/ariSEEnTfPY+EAsSaBYTUMZ1jKo4duvzfLRdjXfY5xCC
u6G35cS9//Xmy52TEt8rKth3OaWGAXpxqz3PuMUly2MBU2SzluFiFDQgl0tWv1lwXfk2SsASJLok
Pr9U5/tgi/e+TsZH9s+qWJQMk0qu15A/lyW9OJqN5N+CSSWxFW26ebqmQgaUnQgsmyZ5E5S4EOgg
SRSoh4xLxKTREOMIl8LK5mIF+DKtei//s5HaqDMEU5A6u3pL6QmH5xfmNmPtcQ4vz15duQRac5VO
Mia0JqR+E46es/LqccgQ9Q/XIVzCncrnPXYdNhBgGLpo4/l1fGLfiEoZR5eSnNhqjdGTqr+YVPMn
SYt+wDg1xHFri3MYM4mu6qJnmBzZqjBeX6pz/gwHcYaW74QrXv2niFQLn6UwIrm3o3iU1QfKOiBK
ZfAWHPY30gMw0SNVMPEjKmcmumr6iYjej/pqBSvTuooihlQDJVzfywQqRY2rJKkjNHNzcYp/B9zz
ykc2CENk9e6eg7Xw961cI4xb34lBjLd8nCrjsKnotLldFS0ofU8CokEPKq1HnO8iqf6u5hNepb1w
Keo51vVAl9dLE0Cn7JhiL6iY9jESVLR3nthPLhxXmiwAePdfwETxmeSb+7pjjhISZepJWWmroe+r
57YmeU73rtT634Yu0b9VvCM1Ee7XOHM4wCnlLCNh6OvhLzVo4/aYSFr2k81B8wwo4ojcxV90daHV
x/L8CEqqRB/ao6bU6aEiSZGYJBw6YLi3Aaf8fCiKy0tjLOLyfBi1tFnH0GcniVv25Gidp539/LvH
VHTFBB17P+iCClMsxZFGXSDfBJ5omJ/4NOftcV2mpnm2nTn6blIw7c6riZsDrm9BLV19/QsOSisv
DSooF2OIMqOG/iQaU1fjKJE6z90ZHapznbFqlPYD5hfo78K71pf8LBXd8QVBAcow09cT8Xpx7mBj
1JMEkVCNKxCcYKh+bej2kOXWW0kEHOSDza4eTeLVbSaAkxFH1udhYNiDgmCYnee1sDVeogdqGoGR
a8T7xTmBwpb9NzneYCiaTR/nW3B3P4X4XuxlExCKzxYYZffBWu+mB4F2PGnL3oQYEarLEdbCDmxv
wEeV/KOR8bxQiV5RU8+tSbSRb9l/wYxdaVA+lmdYaOm7DiAFftxT15eYPsrfO2YVEmSt4WoOIiVl
zWMP704Aqyh+6Uxk2vBV96Bgzmf4aoJBAJ7Z01NilHyzRWqkF1hmFHJXy1qJ5kRnPA+yEzI1C2Sg
QypSKP7cmiPtQlx0KLUGYHz5LWtjI1JME8bRxSYlI52aH5d7q0aPYpmmsZzIRPSogyOKNdxXuTxh
S0deUaq9VNoyMxXxyyXLFCuqIPv0rej8tdgh9hmiDlUck9ZaZZ+L51VhMk7zWd95YdsjR5qk4fDD
y1RIhFbIglTxZRMn7wcd1tUP8VjfTpJxbs3enOdfu6X5SfoROQKIseVg2gUxp2MMZ/8D1ki4F2fY
CDBm6TOcBq9YyPrtsL2TJw7P+8f9PKm6hLh2B8L5nGdWZWn4qUDjQVNsC0S6FJMFU41FgqsG3D6q
eNW5Hgj84I5Gq6BX3MnqlUb4ofK5JXKTXgSd66LHDrZ1XNANcayZKr3fvo5IPYaiBj5Msk+UC+fA
pMWL7uJP78X25UTFN6qgaNPkeZsCbBaUBElN9/gNMXMK2wFOM01gW2SGEw384VWrExKk2hmdBkwH
fet2nR3MCqsFlCWhgJBRFEatjIznlnmCnXS7ZZ3XaNkKNKlevFaBfjsKmnuxq18hVujDJeG1GbhP
prGB4JRSpd+uNJRFZh3cfgNz9a8Ciy42GjBMzh1A2KuJ9iVYemf4pwFGg3H9eoXakqeHtm/v7lao
qpGFkk9LM+26tXokeGttGwPYIK2kQgiE9kDiQhD9nuVFTrpSSRqpIUXvQx7/lywPRNttlFH7NQ/h
GtoXvgdfUq9Q0mG60lyZC+oUZjVIh3MsBQ7A7LGhZvBtGzrSzpW9zwmSD9j6ArflRiPnVSWPYIhf
wRfL7EZzyi8T+sMjCbpV2oiWZX0vLGDDKBUdOXF+uw5QHcn0pWwcb4HRXiyGQ/6nYRAi5XB1x5Mr
uHczMu5Dq4YfpVEZTw+aiYkk/zrYtIbE1m7sNzlV1xiGXqINEsDs+JJmD/G8bv8nINHf2vmjaRnu
dRnSy78mQOpo6ASYbyZVWQ5RuTZTxeKVUtk7J3E0SyrkY7revVGuNn0yKzg/ZjFSC2rFWfZ+wfdv
tU3TcmQ3mC7MYbEwnvTFLjHYs03SR+lPJuYKLEyhB5G4XkA/Ym6FQEdSeJNc5cqSylzsm6SW0B3Y
PkNqihBnO+pXHvS8rCuTfEIAnu8Hwifa2lXYKTeIRfs8zZJ6eUduDQBHsfMYcKqa+cLHoYlr/S00
oOljWCxPMxy3FVzjBZEN9rp7i56G9J98ogQZCxApS/6Da2mLawLFPR/fAQcisyu1BGncsFcmiJxl
xI+4NfOVefHvk6YErnDKiBC55eE/apebZJhNdym9LeCnQAJsLzPWw911Xl5QOg3hPbkXyyNdV0dm
rVLYicoisltA1kNlxVpxmF73Apt/fDHMCKUs4LVt9KCbbOre3/FxzsP9Kl0S9ArLq5KgkTRca7k2
RjCDeAr/GCMsN86EbvLADwChgftFTzfD3PnoqmioCb84h0tTgdUtQyG8JLzm/DFbx/JbzfoV/jRL
QzCNkr1W4V28JEfT7nwr9vtMLxl9XXWDxiqBnnoTB1DUttwbtZrq5RjV+Hc1YPAwS7I8HOzkQNTE
31tIT0B9vqtLyaLMB6dPxkGbDHAF8pPSC1tNkEVuNntQK9kNY6SHMBOEi2RweGtIE8P6Wg/mRrgh
Y5NN8Jr8GaHvdltQ6HIwvCUsqyYlc+6bbswWoWBWYF2CfWcNxBkW0CDk1MlWotc2hBBR9Rj5Ik2L
1m2dKSVV/ICEpVJuQcjQ1/SqbdjAlDyKisF4WBpaL9xRXBRpQjhXk81/bgwA6SYbRlLkdd4MWG/H
OPIoubtfYvKDhbbwRurG0qMFihSKXYtgMtLD+aJzO/CBTt/MVDbEH20Lt7vuX+8C3QBFrXP8qEDe
IGje2+NRSgPdsgQR+QEHX/k8FvgM3PZNGG3vn1IVJFzVOm7Eejo1dnF7emPB/M86GmAexGUuTABJ
zY4Pg467MfjukvKeJUbb6GaShpgeNwqHSYxB7H59LN840uGrMvpq4tZMe7FYg8Wf8LtaKAPNLXk7
uPpUM1QgI0rRcEFWixP96uaeKFMS5RLi74apCcsLerwLf9o8yrEvDGfeZWFW9F82NLRwuR/Z8JpJ
wMcj9tHD6lEcHnNWKN6cuezE5bj6iU+nnABCtv48TuqmKSObp8oP+ju/uB5vO0tfnVSvAtjlax6U
ffj+c/QPfxiV7gbIlzDDXLIxn5pa9v9HoXWPyY//GbEcGJ7khA55w2VeOi630rkDTgo8KbUYxoiD
OPJ7AhH+i/kqcU+78TVykhtjueoIky6XsvQ0hQw0PSBa/AjgAo4s5R2Q2UiKMdh+voF+hfDWJi1Q
Ji/aoo7NPJ5PahEpZeUVHhcfyFuM7GVl/txTKt2K2yOPXkzldCuq1MzrF/5KA3JIh6rMZXgnYz7v
qUw7L0M8IhmaT3hcUe47jApT01RpvPybzM7ad0tUpnV0LvEroSKc1qKp45Fgke7tRFEqnF2DgnKi
gsuhynLP2aNI9jU0BWeem7poRJqXlNgeZUEhkxl5HHdG+XDFrTPr/V1LvGfLLpIhR6iFUsLvkzKL
VnKWj2cfhQr80LpKHX8EDEBY3RDnmKKWZRigtNSU4mbq8ZaQujsFd/LMX2bUU+qoqY8TpWndOW7P
gN8P77Pbl53UR5b51xchsZL1xIxLm8BkRvktnRfz9Dt9fPa7MxNbe6VGGr1Y4E8EhrncmbZi0e2m
NxabCDI5GooLcxS5Kel2VLrCmIYLYdKGOsmXMViXLMU5RgDb61rP6vmsWTtFyV5/WMcQyx9jpCkV
IFzi1IGymrTpH+S6UdBTFZBAEWUky9vOr8VPZKRzhu2ZDJ1OXZ8aOVoskw7QSxPPWvRrU4uhKp7o
3xdAI+1d4NC+PJES6Yy8dbwpfUukEZoUBd9ve3V0WTxnHZDVhJSHoJHQe/v/346KpBreG4XQ15PI
/GGXE8OzNwPnaOgr3V60PsHdWZkanpgVM5VgofVursHzQSEf1M9kk/PR19SFPRJHkq3+SYIrFmp9
eIptmdOaqTEy9+AXobkM2svmVuRthNO5PsMHSgLbsqA3QVrGiTxABor1eRscFbk5qZGMNzmvBpAX
tlZkFimkMqqe+o8z094RNTdM8UatxokQQnlXMHXMJACuFKYhSTz47qf5Stt1GPNaEO8I6nvT0L0U
qSG15f1wfwsBo3m2H/j47HpcBC0riPDO4tDy3fq1x9Ogx7/O3708wv/T//1MWIJ/Az8k8UpNR8Rs
d3H1pR+P1tZE4PMTG5F5C4KwZDLxnsH8HyY2Ow/99CIChYCMyuGSh1OWfcbZoPZVvfMSMFnpnGMt
ko792QVcHstt1mZMvWnWKQwiPMGrFWPyekiSHm6YNnFNJgmYuv7BWMeaMTEUWY+el3dByNTUSKU0
UM/Vq/97O8q2W5nFnubaRh/AFvcWOlWxdxytsc8xT925GbddlD28CFeRpZXZEepz2byBTXGEO1Pf
8kS+EgcMLXHMMJmMktSIubDCsZ/0a+oHg6NbcXEqx52Q4ofJ5fHUULFZTw0/vR4lPSGIFjPSqBNu
zdGI0co1NflzRBumvpMZ9B6pI5Ih8QYduZQVp/ui5oa9MqA9AJovt6QwVsWPhJZc3Eu0ZZk3uXw1
pLwZIsYiF+1Qjnocz/pHwoO8IytwuOr/0QdDruRp/dlwcU2Bzrli4FOux2NUo9lDaH5tcMdj3o0t
QUt/K/Ll4gua0Ekgr0b7aVCZLAxdYwUtsBOb1+2IPHTktq8gTvvCUoOfT0320vdZXa9Ai/GOEriN
U4qCzdpgvj2Ec7Oy+s48dKUQsrXVZRS+CwOjyxgSmIyswC5ub73facLUrowdiVaiAbOQWxtR5e59
obRuhyJ17kPpC7eBbNKgEfxmFekeoHQasd30WToPa4k+9UotP+daQUIe09Aa3c5hvQqywNMSKrcJ
hNSacqkAPuiz+pcplA2U0xuStUpAo42dtGlA6rJEnGM1V2mN/rCaU3QLkhEa/T0f4cQ0g+DbMtlE
zfKKYUmHMKRb9BNAl9BKSEP4ZG8kezegutb6Po+P+5TIyvOTE/Bn+x+irM5PWx9bruFzLTFOmkes
6jTw01jU7iX97th7STUDICD/R3Mm2lE9PLxqIaDYD48skkDuw4XUpqQAPyJsqGMzN0slBHyEnXBR
9HiCPl7pIvY3tYMFdsIzNIFa781/fjDQpKX/74YNcbg9xuB1GACsQu4ryuCQq3Qxz8n31CHcV6ZI
XhkjZl/BmgGEdBcY2Fwf621SPDXvW5c5cHsnwtCakCH9+cXc+0RwvwkBCPOoRxqG5+aYZb8kzJIw
LB9IXrfTaSiH2YTq1v+FdXDM3rVjCfI45Ad83l0kw51RfRNGbcw9CXnn/BZnzEzSOHFHhSMzwK7s
FdCVRaPimH9B+VjEKNDRLyOVkHztQB3VZqAkdqZwA+Mu3tVeIERATfzU/rCoI43ddrJl/d8RW7h3
Nke+QafIVITAjDah3x6TZ9IBt41SltKxKT7Xt7z7QY4e7SilGhkrOtQY4lmrK7ab0Tm1Q0SQ6P/e
EELV/R+bHe4eA7Ouql7w/Z8AbHJuEKu5Ciz+zGrlTh5WGMnLq6okjkyDYsTCOESPC8ijn+hxJM5e
xTKRVFR0Ktg6kwrggTq2MUd7rDs3kV7XkH8epaeL4Yd/VTn0MJc126Lw258UJ2vrLTFWf/S6q6sD
mJ6O/kEghW5be8ksRBNk6j97Py6Qj/dZbTYa2nGDePaEcDeh/WKbynWx7m78mDM8kpH46P2+o/jN
3r2R/jN9Q0BEb8IlYkA1RmC//5coOd6+M8HbLR0/TueKBc2V8Gz75M9j4jHlqoFMV7OsLYYLjIRG
IRzf8hdP7+t9fJsNdAHfqg6tD/YEzCrU1Vb5AKEHlj+XSYuD+Ao0pPNhZS1WMXySjQkeYksMTDeR
gggc9y+6DD+E/2wxRvlmxzbMzuwEBxOw5HhmOomSzScVtk1UKG0+3PDnxwYZQJxRKDK/3Hjgb01f
hnahGM5AyDWIO6ykbHQsOlkd5zpEH0ap8q7XkYLpDOfc3NfCRqiyPYOHflt/sm95RzHwRGpgcqnS
qPBfiBFr3y6B2yvgLR7dhT1w+mE0E//y0pRoDyIyGHg47ijQSVlN21lDhdexQz4lKn2/ABX607N+
582Qg9l/B6FdDZVw9Y4WaC8GUnVx8dRqGmA/FaO9+iazgvKfNu0XbhRD/ZUxPobNdkB+cbtLxQKm
FDQghh5wjx47SJmNZ1UNjXDA69wTv+sa2Rn89IgRNav8VGxVsajTT9l2VCH9gByKipFbceSYIy9r
L7US7LnaHaXxBrZeyAgmtgzSEUBVEcQQBkRQ8z7Z7rZpQfhp3mWuqY6XafpzVnJmzThZL2eXtfOo
mdzgX6f8kj2pOsUkacQALGaLGDupfbcHxtHwWRt5LyHVuq2Tfijvl+9l3BFxOb0TSOXW970g9Jmv
/zhKrZd8VqgcbIgo8UTpMa3JzQEnU00pt2C7hmjMY54Y9u4lueR/QktfUv2ERNVA8xIf4j8bIJo4
8aRNcup8XhvEzNuexj3fDkgGj6JFwBgBwDtzqxsQij/K5Ke1Q1r93LVxk76CeTpgv4tRpcnkD3qh
txi2U50jF16vfyX+hGjg2giuFoJmUyjBJOMPwqxT0+zn9s96lWVTSBtKoCwJHeEzC6eaRh0pwgij
mmi1cQ+K/cmbxoDx/jAbNYUC2DMebeAZiUoseWlZ1t6CvQhbYlbawBEfr9EvosR1lpwYBmP7wXb1
TK2wNdAWdOeKAwlS/8ZwFHQsWcPMMmUK1M6PnxVCUD9HodqIodufm+3A/AsxI5+hWsn5jRJPYqJy
bxnlRoc5GtcSehTSDCKuCQHh6sEprLOzi3Q9Mhtl9fzZXmExyfAG2ugsV+glTRfcQPfL+7vsyqh0
3KCuTCcaaeJynk8KDejATpbZjc4rIi+WTznIntpAsHcDscaLiwjTqOjVZXPqQte8tB/kpM/5GxUQ
3uOWn0U7KliKdaiTU74ZAet33xkpAvQLAk5RF1UYlfC9m+3cu96PTGYRZLgW09xEsDy4CwqHLPZJ
hqEBVt5UkLvCDvdBOwLYnfykPxhoHCDW2bSBs6N7PqQl8wLItbWwmCy4FVRn3eheTPXtCPq+YH3n
09TreNaf/tPK1/tMM1QBvbmh/i6FzY6Wpm8+ggHawUQ9YxmuK0rpn0PnNV2YQI80tlgskn+kq07e
X93ijax9nt8u4uvF346/iwVL4O19iAEchsRQrJZGl0ntn2FmtS64+O0yS3/J6J8T+3+G9TH34Hdi
/MUk/so69j/7UOG0SwXR9UDf5kuuBt6+NYaTtUjq81ANDAR/Wc4kvjPqSiCZ+TE8Uj11aK4t2s5d
9kOIU8JsJpE3+Cu7mkS8lLWEdroYbaXo4AoYm+w3my240WTTZPdTAAE94CMUiAV7PXPFbaAtMdoe
mpCnb64TvwHpmt2FrXiEBhuyP3Q930mnpRSiEWsckMu24V0dtyZPYBo3ZdMrCYU/7Lca4b/qeEt3
L+857Lo9d15tAIuI7xEQJXuWPZ4V6cSgcsZteBY7CrJ8myMLlKI4sizFG4oSY6baBDnDwzkQAISI
mMYxxtSmWFJBCporCXzpSpAo960uwygtVdywFQtdKbVLINx6z1WqgjVTF5AfOp8AbYabDTU8ObkR
/qE1u6C9S8amutpK+ra7Qhhvzt4I9dlIWBwpnAIzd6d37EWzYXSRth71cAsmEzuXfB5Vu6JNVDun
AXN40p45iiMce1ekboyRR38jvosfAda7yfT1HFx8fYxwrNiJkFHv/FKxZighaMXBLtco3mhM3Jf+
lwrw/FNXiOczKPqwxnY4C3FBHtZEHnkFBiND1ICdpvYETYMdTtO3qD7bTcJuE8THCQ3w4smd/I+s
z6jh8yXM1se4USLJXY2CmJBmBhrCNkvSlnbiWbJatH/t0NFtIhR8NAj82zz3XOsAxVI/np2/fFHp
G8vDzElgpkBgm26GbH7+b00DvVf2J6gZdr+Mu9H7wfEMgESTYA0U8UZ7/sC+LpWLIrtr1fxNcVDR
BliriJ6fXCTl9eJ43LEj86XhzS3sZG+tQXpNnwyx1Jv5mvngby52b5TCuvqJa4vENLYkcdSdEjgP
mvX2J6w2TKrQnulXMz17dy5WIaQxv67+DQkW2e/RjsoIAlSDa6lNjDdWE+0MSqMXopRP7Xw+/5Zg
eCuLiemwsyZYKHbLwF7NAo12+u7wjmm5ZNAu9WE/InpW+iDcAyXbRaykuUA6ftcLPCgZn2a0IQUN
KgGhJ8kQWJUu8FxattzTvKDn2tFjcRCKiaog0HKXQaaWxiCsYS/zTExGwmEOJITq06PaZnzhZT39
UdG7kh+e2RQAJiveg5Q6yrcKZiJrEiC/csrnlLyiBjxXBIyE83fVB5tO1a4HF4f8L4HC8TEvJ2E8
hU/u7LO6Z7taYVniyw4niAsoWvGj1WksAPi/1OAIPqjEWJ+iJpv5UrPtH0IlkbVYW8tyr1Hc2WcA
yGDFl5avBGO1HUOTJZavKdB1qDyKC6JBUkO8PJnZWvGMYv/2V63lKz+FOxX4NrCXiFXxoWKb3LjG
HugoMVSZVQf0SwyzFSOlp4TU5qdAFC/z7vcv8ednzSG5NlxK3Ry+z1twOjq5FAYD9oPAI7J5MZHe
/iVzKxcShXSbjtjVYY1TMd81X1POXhPGc29dpwyB8779ScUglKcdA8IjKdOLJ6BoejbmuLXJspiz
J4zhYpG4tQVl4ra9EaBytbXNbrNChyXak/miTxrljzzvqugS2L21m04s9g0Tnt7wAdcKmBMb2zI0
18OwZlcr4+OhZM2motyT7gM9OixXtlcKm27/AWDkqIBD4eEnhassQu6a9N/2RJFIjHufSaPHJ/H7
iTwOKImdLK1HIVlzdestteSOtvyhPhhP03CGTvCsTRuZR41uYHVk/pn1xrsHqlPchY5UhhK5esFe
IZql99FQoseaxtDQH0nCYcuwE2k7WepPw/rNAidqBMVljwsVHPMOSBemEfEog+gz8ICOJS/g0b1Q
cPFf/GMowsYVutom+zU5SYsD63DDb0a/o98mQTCj3/1TTKAvBrc1lr9mRMSYSdlHzNjwSg2Q39mZ
q5k0cLQGwqvHt12nIUbw+nwS7O+X2Dz41QvjZES9TA/V1Lj5LLdBZS5vWNTRD1z65iVewvRm6BzG
AVi3l6Gh8NWwFhqlaxfOlJhQBg842XPTo7CoRKS5V54bzUvTM8y70QN0fBh0+UtARs7/4EtX7A8J
/kwlKoQ70z/VzWu7Mfgv90m+eVYG534DwkztX9e6JOCNm7ODsI6IIXCvwwsUIK2HXszEtwVoYgmK
6gggmebifcrXlhntjheTJSHEM/hzJpv6Ia8O65UlGMAIKD+7ZkdDyg6v65X29Mt7NJSXx/phyUel
AGOHMXZayIATEVN1iWZ+G2FDPbUkAzP4DgRPbIOdyDHtVSFJWyei1QUu8Yle1f3qM7ZIUFaCVMhI
b2Q+IqUGystRizs6KsV6IgqSZLFJQqXp5AwDyxIQdILRNf/+b+cu77lArSWnC5BTYyYvLSJxgbBY
W9bn1Ty31k3Q0tUMO34zxCd1MhUs6ylBWByXCwy90OkUHNzgDp1nEU+zPq8rF/wMLsV2g2kZkFWP
fEXDW/alpuA3witHRZQQAMo3gBvGjRGmFEVJZNKr6yCW8V1UmKBIrc9y7KJerO1gLF0d80oWj1nv
JGZ5hX0D8/iGqHulbdSTJClwj/7kPdegFSfbJkuIRKnY3WcNX16XTiRy+Dl9Z4GLNrEqubWtgY6A
yIvhX8dj5VY7pqzk9D1H0YUB3dgB23KA3oY8FrCDdtnHzeUQqc1OOeIc0BwOEIA0tWiFkPK6tPyY
AK9Uj1+UXy7wIkFzD7u2kpcJDA0o0wrdTKeK735mQ9lgO3IkOdkm+z9uiQBlgT6yPcm/i8uQ2bLq
TBPziXWWHMJKtbhjiJYz/qu4HEez6KFHP/d0L5vBcB6H9iZvXig+CJ3To+ofZ0y3JmyiaIHtt74S
/7nWYFiyrPPMSommApyhNM+K6vpEmvEIu8u3aVemLeuVvyG+icZOzuLD7Jk8GLDCsywsMUdIwp+P
F1J3JlxYsmVyI4bl8SvHlJdhmrQN0pL4xvmmgLDtUoCg9ZUyK/wsBq7Dpy+LA7/EUcpL+6DWUQpb
JVLEfkbo9OPP+mJ94mkIGZD1ONBb43knYT1A4USt1W/Ok6FTc0sidJwsN/e8JluRxmQGXxxK/Xql
mBuulzDE1Wv+5HmVoVmgdbx+yus7/8W4c5eEDix7vagyslSdjn/r4HD1eTrXcuYC1JAaK2kVE5+R
VImFmU0HJk0gG3PbpZn+w2aADajpy/koNxbtckDIA6pBXERTnUIytL9L18N4GMnHF+swexhd8uXI
dmkDjocRnhWwBLEzEjBXKWxH/ZkFAdjg/ngMw07T3kH5ACUC0/pYtkwKS6i5LM+FT7XccNs+XHJC
oBXe2K38h2MspJvviMMHYiLjrdqFS9U0o4FIRnRKiS4Z23K8B9zHzl4dkwXze2umAYplHMDn5j6y
D67X10OZnb0bATKzB9tV9AOADADzuHmzvsEz97izHeMBWIug0OLPea7d/EGNDDDbcfTuziFkkOB3
LE2t2StSeHRl2wfqlvk8ZgxFfv7ZWb1dveaqGzfq5YCK4GKo+obZPnYwOthy9L8aHDsoNdBZeVyW
kIHVLxj/AbD6uWfRPS6Tse9FmYjOI+1strVoJcmu1t8uN6QDDgKAbMWSNXiPO2qz/LFLBbloW0Je
8zN6h0cVP97snSopUCI5aAr4LqTQ66SzNI/kSg7RHf/3v0XwO5XCNNWn97xgHiT1pgN82yDEdQ4H
M+yes+Gfyt6UYdSeZx+fSc1PqHF305Ea0ZHhal4kpAoA3wFKys7owvarpjZJqktlmxdliT4T27dX
vk4hXqwvxXA46pVtGsexyvh0mLSHvoN+EoPYmerBvnLJo1A2ybHKL2UOTBcxUNnXIjAlsIqlKBC0
8ge2XpytdLAnP4X2VTHVWRO2NRBdZZ8qFKeXLhiIlrFGZaw5yrcCfTZOZZ+AUO7Uo5gimQdGqLnA
NkMhEKXBAX1s4gogbjrpkAVVergTFCpmzjEi+adD/Gt/RxztVfCeUGRxWXFwep+SUicy8O8GYTSq
n5H2vl4BzYX58Wh3OpKK0ecyZ7hGrkmG5+EMigzFY93el9f/qrQOg6c7ubSxYpls/zC7Pub5GagM
6m7czlVgK9E1bC/2THK1IcpP+CRFfSAapTkGgedelYQD4ipsa4W1bEp33f+z5adPSyfc17/S4BkQ
CNy/c2Dat9V69JqORrQ5Cc7M60h8dqYsT5MtbDJlgsn7jShZEeu5r+pQ10n0vZJWMzMYuewAeafo
Lnq2AXDXh5MvpgxqKh3/McqlE8R5aWPskfYn0iOspHIH0eQBffsxWb4MeTuESFDnZZwYTChHC5Dc
Px1NvVyWBr6Yr93H0A0tNVEAb216L6MPPKF/4C5IRYfsgwAKpg5+GAATLousGkjeMbDtlTzJ7FVP
tkoaHSSBFSpk3b6wO0x6X5ygya9T6BA7MaJicUXa8nCynOQxwO5lf+9n0w0s2tcs6t5xNzQruc6n
ZiEGUKVE5X+VElz1/L4npTf4mmxgKu4v/0Iba3fXaYjmyn/8N98ALuYAvyawyK+K7bCIqjti1MjC
dLAPPien1C/Ea3xrdsX7kigbGltbcQo/1tuZhNXj+nH1oEussuTkiZxk61riVc2fcGozjFdDdEoR
IRcgUfttpL9XhWDXT5OMw7bOCxfA27Os4ajAeVhqntOmGoDzNh6Zg0hEoSV5TE9iTccJYmpg76F+
XCiK7K5e2PRLN7HYtE6uyFY7G00p/ssYE1NNK9ao/9Zi0CwFFalC/Xn9pYhi3jv/R2zskoivQuLh
KSIwX6Shv6nM0+k7guX7Q+LOKSiEwpFMJVVWOUl5OLkOCmRm+yU2cBnk4MkduYKJeQr0xgAFHvDG
QhcFg1EYPoPNbBhNvcJbDJx/k8PZQiX0b5StkmJpUH/24o3oZuCECUBLFjW8dA3V2W9gNaJZmuFv
YPTqZQBlHPhWIx7YfKeNZBjwSbYBlzJSghu6HD2gFsMizTGOtUVvTxPmeSEMkpenlKFjzmZKGOem
+Y+PvMfLA/wxdlXC2kSjKbs2pOX3gV9bk1mgNzwvoDgpn3mjs4kyM5Wn0W1+zKIZv4aZT7E2WNGz
cfE/U/QQvPWM/y4imOzaWlfzdkjgxV48AuEN7pZd+M3Pbn6gQIFlxdFce2PlcZT0X33KXqr8v6Hy
IVsUmhv8+peEZsAlfHS4vQWeUInH0OPxbJg+5Ya3850BQD18MQ7vbWznusGQp0UMHjmSJRxlJPPa
RWVTR9vIXO99W1WK7MBamHBCj5g0RwO+N3E2+jESxfNxteu5oNgZ+yEoiDuFQpP8ytF5uDV0Mmg2
PdhbG62KJ8Po2hCxbkUwBS03OIjXBYwulzrZ0rojm7zlnEH7eVgAW9/scY8rlKIYXN/GFIgG+xdf
HtiuJJqPSDBmkqkOMtqAxjxiwoL+b0o8+a45PEfh/3jkd1t2Geq/0P7nLh6OTAfpJUpGeo5twc1t
ZaypIj4KfLb+zQkfPTazOOrLjnq0YSRen/T/A8AxHNofSoXWlgPo6SC4+B3PPGOsYHDeLt9Imzy0
Y55Qwre8T+EmsNT5ICc3Twkg+dnbzWEi6Sap/uToC7zk/K7Ue091k4+Z/VVgqp5YYUN1/cU9LLth
1ot6GRiTMlzu1yZg9y1pZNfp4gXK1TOUBVYip8tCnPJ3vpUdM5MrUau1wk2ldUiveFNJdL0MHrwc
1JCW+po34/NT5OiP9N0T5bZxH/BD9wMZfaL9L8s+WgFG4HvaNrNQ8jKoyrgeEvrVwyPG3uEgBkRn
Rf3IqAegIlcsFR01eqnmq6q4655xQFJcIERiWJogKuYxR6osvy84zBF3YWrL4AHiEOcdETRwfvfS
SvFgrfvvMleswjGyx7tqG2ILInqLWQNtkW+N3oYrgROeUkOIua0sWEfJyjwmnZqz10WOcXOY50xv
LLbdC/bhHlYD/cDCaUq/R8lhwgEJWpWPYm4aOwgFbZ6KGy5cLVnX2SbXMWpyGb8rYSKk463HEQLS
qhhvgnYU366PjiQKk4aJ8r8KS3A+Wt1QgO4mZ80Rp5hPs9aUrhnmR5cNGJGzXu0qa1Y3cgabnbnp
2fr/vYXhiTe9XmZuJArRy8ttOvHmx2BHLjdy1MOhAVBL7JRHuHY2Cx2DVPK9zqOLtE0KZguSwwgr
fECw5AcyjnUc8H7CGY+ytD9Qc2TtXzl1JwlVMBTYePFo7XVG9poODFh2ZP//WUb1/g2iCxiwe7Fv
iJDuAjEHhCld5Jd2zmFTmLWB3ZkdfeXTLypGyyh/e9x8mzItnRria+jqxNsQ6fh2UoEMqiOAhdpp
70SiUOFwiyfynVDRQb5XFdHwYrSO67s9iWyU4C0ueky/DqHsQtQBpWiMOLej7G+zV/hcU/vuZ+Wf
fNg8CZStLmIU3it6/SVX2xBG6xJQRleymjn1FWZdXW6HO9JsjikwqlSJXGmE0GuTMk+aW2QzRdIz
w4atC8+QR5y3bR6eeda2w83bF9AUS5j1wraHoVN4K41Gql5SdZyyLVvTq8MDcOU9wBlWM4FS1OQI
b62UwNULkaHjx5rLHr7O6l2b4aIqlRSf8K4SgCmHc/7zQsxj3In8GdfM1WudWhSvRhVkVe0naClJ
J0bTpjB+DsWRCSMVWIDVQghpvwYJHXe/E92UuaGWFYZOMqwZQTkdRDVpARhu1eJ+5tjh9t6FWd+H
y9QIiTm7JwS0gsN4ZkEr7HBxLeOPHs2jjVTzhqGPzPAYpl4R0/xw611vOGlE6o4YWSxlkoMlNXWn
ZH2URrt1cSZAV7oJld4CFVrppswUKfzhGtALOZSPuh03Jb8TRFyARc/P+kxG0vdLN0eXEDu8oqQd
VzzNL01c4hDexxXH8G+8Kexkox1NRiOAVD2G3j+4qVhbH/tBzMDi84NX4NAtMBl/dbaa5dqh4sID
eNpI8AjaNi4lbZyUPDIIeGSkTKCg+3jJZoo/O9f96K7vsAEBKQi17ongKp6haCIVnak0c/616yww
SRpmtQ9o3k8pLDT/NjWNpeBSZaJq107USc3yQl+Ej33I5xgGOpdZur2fV7nAosMZjUw0gdEz17RX
fjqVTCAF13N+bvv4h43w90Ez59/GPiG4XdVH5S2LMNwHhFFFj/A8iFiLJDgDHO3iJOQGr7QbeDGi
nJbj4i58UE0RCe/WD3iGAUPKpM+qOfTyyuela5DmESYnmGmXV/Hqzakf5GkuZgjrGyFJGPcRxX9I
DZ2vOrrZHcxhaKWgogf83Cmvg8rt46c/0Gdc5w61nzmd9CFkMlgRopPVkLFDnahYNKgQwpWTjBH3
seNnFFa4HJz2tcVtDcWZXUN4WVl8Tsf6sxVmPQ74ssvxUQKHzLX3ZiBcW2eAN9XRnXWVugXcMEwf
XQSSYYHV1GvuqfOiSm0SUGIP/iJUxStjDQUiPpqxayPGj6SaAPNLd+aWzct1pRRxwgpZvuLWa0fY
2SkjHopTxWCQkzaAO4G4vYueFC/1+b3aUJ3hwuRrL4FdHoCEdiU07izcvCVzxApqDwigjT/J8odW
oyImJ8aFusEH4+laGf59mAkI854qym+h6z4ds84ME9Mu7+TzibfGhsWiuYPk4Gl2Tk4w/xiLia7z
xm1nJoGRkRobfy99qnu2qqLrLiefgX+wlqeOR1pAqArlkzKF14VJ6khZVCGXdgqRCUGc0tp8IAr9
LwbJ5jC2s8Ihb1DGyjr5sYW8HzhzRd2p8LYY7+jvJzmTh4JXDAlFI2KgoUYvc0MSJgnFzx+99zIo
njXFJSXdWAYq11jWsNanhupvSb7XmsytJ6aHfnHWmpfgA9ZaWTRnrgekc9oTclQssagpTUJ2fm16
rYE3sZScEsycDfvlN+1yuzU+L/FYFy9TZTWt/UGxzBfzZCKPLDLPySmms+Jrc/tfzaxSy9LC633G
y2JUEFicYqAU7ZZYcZnupOiKGdHu+/WmmBtMDpX9nHT50/pTLZp6hOuB5ZE1hh7ovuJ4zySv6Nmd
5bnRbvckL6gbVaRMCAz3C8lSy/K8VCmvx23sT45dvJGd02NokQk/WWuMrjSeMd2kt31H+LL1ZkG3
DmOkn86DP+M/FRVOEJacv48f5lXJSs2D3QW0NGJ+p5bdfWRLSDiyq2FsfIbGfJYSzX7ZPwvRl522
NeJsQC1bDxSglyJQGCTx+jfqAt6uvooPddDUaZ/p3BQLPO9vO8yhV8OBP518/VyzQBJsikUGgLqy
FW0tioXLD9RKiA5pALIhKkwVIXubA1KdViJkiH2+FNC6RLWrXjP9nz9iEihJGiYc8TjRGrNzZlAY
dWjDra1rlOT2zPPJccsl77tUICUe5T1E6y4U5cMGY7CNrgfiTbbXnygpX9QCiUDm0+EKjwFN/BMQ
xN3kev7YAB+/aa89fem24MLyG2qT6Kr9cW+dmh8rlPXksPxvp2brcLMUsze/Du0sBaoaa5kHicGr
+iZOJSrER1DjLUHcRxZoJYVkQzYVDOA0B2Gg/mRsi04rgPE/+8Y5mgmHVqsPuRfs8dJz+jX5J5Oh
8cVMqqO4MLDyaxvDhuZKnG3bMZltzAGavNYEablirda9YVW+zDpWRGIcVUkn/D+TJ7+Li+vK6kff
jo5iJ52LYgFY/0OfknD7ZkZwLZ7MtxgVUVnUJi+trrqGWNaU/tfEFGBBlbPBgOGHgfQ4Oo1rfo98
nyUUxbdclrVa0qQgXdxUVxf1z7PIcLtQoDcODjN2prSkuw6ZBQfRbwu/M05V51LyWkWaMEtAqWZm
Lo2VhsHlwaoSAJKcV24fuOP2LGERuNpBPOqTrD7ogs7OAMZGEjtninsRmPfaH8DFqb83+1Qhkyzk
+FrfGU5j6rQIPnOh8bTb/LScixTcgP5RQwSQRG6BXIfkB5aFt0qyxQs9FfX/5ni4udTPDMZ1ycck
wKghUXt2HFlP3gH7Ry4xgs1TRC1vs0UeHRtWCs+3tRhlS7GPtgOhasaOzBSpBC+03nNI/sYHJodj
7FORio6/IfXIYC24zvVbSzzwHpFZK7fuYiZ4pI+iOuO3h/KlArOJS+ZkbXgrAS68zmpVv/djhsrp
AtqMX153botA8xQlf3hMAXBht8G8b5IFNdpjVOJq/enNux5P0DgMh/kkC7gaq5Re3FPorp/J66WH
oZ96DrTdDrLyWy3UzYaM4HtcRIRWMOom+6Ubn8Hjsu5i3TN15uyhPOl7R33dBrlVzyBVYo2QMmhS
IYbHlF9W2lFvhmQl4M168dqDCMOX7r8oflXortfnbDbZBQLWyAatDXGt7ghnWuAgYR3h4VrWmP3+
alquuekLaGljPy9jtmbodB1uWF2ikjFpddGCpvgNdhXSh0+CvvXrtilzhLnELb4Q79Jv1ROfpooL
AD9DF/PoxPmWmkd2/520/FQTXLmkLOJjyZr3ABuaBAwLd+K1Fe/NUuIp7clsTbVYRiu7n/KwDFJy
Up/5oC2slQU14l4Ry5UsRj6yV/pzHkK4qTbC8By9RtGyKr0+naYiG1CvMxCj1PlSewJHYPn/RAmT
M8j6ipYFdTd1tNZEKffDaLz9292ySKGgHqTSeL7ZtCb0m6naa0TgEufpdr7v+RG5bIrYZmbPIx1z
QgqF+03wkFdRY/qie4zCl40p4VyWTQdzYeFJWGsym5GLTqU0lTCVp5JVt7WcwRSHtIu59xaPNtIP
HXQt5rydjQWii/qJIufzudZ20LcwZ3Iwv0J04gdG6WTs1z3SoLhEnfrlFxxC9aHwHQxchcKB4ly+
gfFJAZkkDW6Co/HGx2nOKwxJqEvKlS4Abhi4zvOlQCheTOqUgpwMH0IW2znjgUSNTXXUwut9wW5x
z9aT2UMa7O0h+BJZCaOnZhV3z2j7xChi2JUNbngZzmOmLc6sYVSfk0R5IoLnPKkd/omQtVFKG6Jk
/9I7ubzAT+QuQu0owvz0JNr/ntnLwjulrlV1rOKf+t11SLv8a8atVz1MJTcPmVlqQXqLv1hEwjrz
rpzeHK+rhKTIF7xK2ekz8TspDzV/0bxe84VdADAcL4cBYDsEKH7X7kO4/W5vSzZCmr+fL8SRmwSK
5RxKeBTcNQRPzKxVCxJQgTBbb5pTqYj4xHfUQSv8MWkUhmjM/i2yGVDdM3ntZPCQEgWpPul8nzCJ
CcoAYXnD4qHLlrNxapA1kJpyqtViUuK6BXa3t7TtAvQ7tK8gTaDGsViy8Ng01UR/Zn8T/iAbMLVM
7IzIWqx6cTPtIy04at7hrMvqNVy5TyfwEmsuc/hIattx8prPAp1GBrwWfz6cdGOdT3kOPSJrTXqd
5sJ4PSMgo0Nw/Mw+ervsCC5X3LXXHLHNhxACmRxbX8OHm3JgY7ycz3xg70HVI3b8akKAN0cdyQAd
2G3Kn+AHx68WtJGp0kaYxRlOTD3uD10+MMxACZOjKxcbijK4p5rEcC3a7U4XC5KaOAFJJQxTqxLq
xG/qu1kTe8+WXTHYFnNdcjDtdQ6p4MWaBvo7qe9JJvAGWGvSUHKklNhBgB20Ac7Bbp55XsJSais8
TBELwDZG3VItAtLkL907vXvK+c1jepnDZwRDSmC8B6UKD+0L9mlyUFqf3Th7bQKgr+BaRS7PPX2L
uwJSkxVkbIoYuUMC7LB/f+B/CfGX4DQnTKOAW4q+zX0m9qt0aUqhZrNAxknIH9FaxVChH6jjdCBP
QfCdFhiLN5MhLzsR3YdmHUc9eS1X3/0EBPkV3JvR7Ju8cIZ/E/uVT0Nvg5Gm/UhvqZ4c3Fq8/GKP
G1NkRaH8w6l4LJEvGYyt79lmLV995OmJkFATswB/UyIyXyeNPZMmF09Oc9MkTli5TEZWrjq3kQMp
zFHsGd8dFPOM6+z2mwTH4AGIk45Df1lgvpx2UJxlv/R79Ns0FdGoMh7952omAhEiNwKVsRfTiVGy
Ptq1ShF5iWdjpxZHvw6AnNClm328H1N2gf1pMpA83sTL/JNT23Gt5eMh4UD8Vl5vDCjpwGSk8oNK
2FAVYTQtMTdww+3kFqYQTMegbfNdG6Xn2T4aH1Vi3UMeUkn82lyUCHjv62cZGY3S57YwOr3/QSLV
T6/seZ5G5JYohutnJej8cG7TCnbM5Kaz6lK2Xe1wShoCuuz0Vkd7v2J5BLXZ912YU3Rhui9Am49r
N9uxNryM/s+TmQvXywFfP3qoJSxw0qpXNK4wn8rtDJxRoVYSz4pM2PvwoQ1eSVjbg+wZqG1AO1m2
r+GrNwl0kzZp1tWFkpN0c4F620EwEjpr0fKjvMt3JRELhp/W/B2RlhUCLH0U6UuHTj1IFgxAJSdL
CJc4qmmZYpKzQXcqzJ5xAWtnLsYZLRAcUhVVi6OWvTR4vWyPXiF0P1CfrBHaCkFdT5ma7Ckcx6xw
CRthNGc9Ph9xSbTpUlABfAoEtG8e62EUX+6sigvcd7sW+h5VlDMg5JO61qoBPWMR/RKHFU8/HoEc
KHvuWVW+pXFI9Er2/K+zjuTJ/hQpOIS6jf/fG+AX1Eyn1v3TtmE+veqCQEy4c9+E5/eYcGPxKakz
/iCymGp/gFll3YKNknvJrVzdZlz597Ve1nW6veEFp+kijNafabEm6+tosXubBtv00u62A9kODzFV
xZn6kjQ3e7GYfb6pzjjFUkqTB0M5nA8u0K7ILfRq9OQihApJd3Tksj7a9XR4rF6oAALtWif5peSk
X3HrZMjfBpzNUUK+WTwKzNyYh+gp7TzoZOeOaQns6KGh5gouGo+u6JoRCe8PRz2/40kFckcQqg3u
Ltbo5pNhnAYptJdw5HGOjxYAcb1cZ89LrSvFXNRLOIpEy0soCBOVLlHwGupHAXG9+PiNI38/Gjsd
7vempN3I0qO/OLuCRBEi9ADxHABBoBtKq2JLoukXeBr107iR1FMGOv2FBFmwpAwDN+3Mpn3TIFBy
iNq2kxdMWMfE8TQEfU3Yh+YWOZwE+9NEPTi2IZyYdzBgguk9WX0Gj+pNdP0febBSUr/pyufteC3N
x43JZtcv5UKKWq42lVdpPuCB9HcjJSO6dz8lM4QqyABZBz8ZwYZlN0nkpILgpxgCyr7JLqHBfQij
RgSnJe3mX0Ip/buHzWCIIUXOgI4fcI6SOrmgkB5oYUrgc4HS1zt1aHuQfMy0SMCa29ByTycx727j
XrW0pfFTqnVJgp/NWYZNE3pdVh0Xw9P+lQf2hGCzTOQh0gg9uKZYsViAvwgdsTZDEZtHbL4YK6Ls
/WZz2cxTvQO64cagF0IzivAODBK3f4SjWoeaZxAtGizpmYpoTqd5VHxmyWvAZ+5FcdaPO+6TWwJn
ZzwwgGsZXjmE536yvGKiWdN0Mfw6VUMPUlgYFYZKkY451QWRoMTaiqi5hMH5rsF+xRUxT4LFZ4dY
cXwYms3UFQcSNNh1n5vasLp2dGMB6iW+yf6yRjBDOBEw6udic/M+Qg3FfQoraXvIk9stoXGv6mhN
cjzHOmMIqPrgwgcVo+SL4PQxNQmAnt/vYfuiNnWQh10rpF2aUbLZ1UFHs6YYzLrcdrK24mNsU8sl
le6OHFgf4CEg4W142Tncts1RMTnnM0dGmU8tnxLZUcAkogc9R2Zi5Lam6NCGAC9BmwO5Th0/oR/k
azjdCRBp4a4iS+W/5EH1hIW7Mt+NpGBp35/bvnOpkBURxt9L1kGAtr/P0P4PdW1vY5SqoDp8NbqK
cpep3Uis47dafYE5SrXgy3WaWBQVLKorrDnb1RG1Ej1dnQscONPZsJbzQWXJTlV+ZMVJvKy4xDlD
HxoJeMhg6usV00WIztB+EOCKpEa8zIh1F/gVTdBn+Wz/mcULDgQHdJWP5s8LhkWv47bX2QRl02bL
A3PD7EIB1jkS+U7VhFRb8kHIBbR56bDj6LzTGhyKBC8fUMfFVe/wpRTl4DPN+n30Dg2GdqdRk+bm
54o380D6pFCzi1WgsdpEcO/QWe12fpr80AyfdIg0K++P6hFHq70kXzl98N5S+5HuV+YmsAG8A2nv
LfOJa/UbD2XgF4qZiaSsbwRN8iTEwARRn9OpA+soVXet6ahmqOl/IADLxOT7dEpo90ijMrXxProO
6gJA//PaBqlczKzl777dxX+uiGjAau8lC/W2UR+0NtEdhKc1XbNNF8ollaPVOGl3UMbKAx/C2m/P
8pUSEOYUh2dX22I9rBmh/ITPgg5WG+snaBzW/MTwrXksBiwFlpsSCUIURtZUzwQlLgqP7cD1HE+M
BjM8FXkE4/pTrCNwstgeIZ8I214bJyRAHjltzOMFy3mVuTkGNvuPAb/ylhrzLGzcy8usKsLWygq/
sxAY0hN8DDoc2tlA2WB44dsCfW5FZ+nOAq7ZV41w55Hqk5rZSu+bMtMm0i2vnooDGWg/ZdFlBQVN
qUfoXTAwwi5Y/yc/OyrVbhl6UOlrsLe9zA4Jrwsuny+e/v739sGodb1w5MuOi59OTKcWpCfrIJui
LxiYDGM9qSFPg934JbMTgJtpW4NuZhmpLmi9HXIv7cllZg9znbcm18nHMBbso895H1jPRwgVTP0j
IoJXdHKYVrwxuWeIG0fOWbDapyKh/+Nc5sDIl8q/614jHQbfCnpssqpX2jLAVkgKMR4jr7GqkUxf
s8ZmvJpXuULLmWGy4ZX3mhzVh+8rhbf+juUBPP9MsMmWjSziAmXVa3gFTRc/vk/8xoJeQF1RE7I8
VGuRt1GbdxCax9podc/q0YJAeaTueRxoCCpaLY2RcRxcGwHsbmQgngl6+4fAP+VkU5FTYC+/3TAB
abeDKbewP62yxBSitkqhWn/5P6P+D7Yy1Chif7jUI5dvyV+LIgJG7EZ8lc3zZP6oftAiW/t1apGE
rwtr90z7SET3c3QHAtx+ePXiBjHUbNzbzZXtohkVEyooAJfdk3W2s44k5e6MUDo4x6zRyv2ApPHk
37oPkspaDjFSbCgZR5O4BEm2zJVCPsGJWE7HVOoIugErAjzZHeuxNN0yHg3bDW04k4hI4tzOK6cY
4qbtoYhGG+cYjOHhGzaxzxI4HzLJRsPB7sHeUektfibd+3I7yxF1k/ZpUc8Gse9mM2yEMpmiR428
IeICGZvaAlvNAn1+aIiuuwu01h4nsaRZm5cHLmC4cpbo2xy5tgEVCkboXQQ6/bR2le2wKhv7G5g/
RZrfyUUrUdGgHDaXECBXRBFLDDSTchdnF5nvin8dv2AS3XMfUekuSqoEeGqS72tUOp7Jd6YLs2Yt
VRTwoZGS5tt3yqvd+WQudiKcNpFHPWT/YqB1jUrKbrX21Qn7kvOn6G1IaNK3fEGZ1Bjyad2UZgeD
vwAKjcRlHe5X+yAhpUK/EcOg00tADSLrx8lC89KoF9ptbliGjDMKKXQlfU8ZXzUni5OwAgN7kCVx
c+Z0RqnaMVaVIXHsd3sSTZhjGhawSAkt/LxpDRmD52jwP9tD9HrdETrE8LYXxqSpjQhBjulttD4J
Fj29spO+KLBH99bwFgDfKQ73wwLP3F7HgxaUH9lSAA/1Jq+We+u3TPfFVqTHLdMqUsS9+HVK4sMo
MdkSZUuZOH767zTzyQ84GSwB+16HpRU42LyFlPn9mUMId76QrlQu6dTDf1DFMmEgVYV0XVFYcZcq
DvBcvSr4etmuKlh2uMLsljE9HSQOHJTo7z7RTv31Qh75HAIXWN04vN3ZAlieO42zFkU3VjDdLuR5
w0JVQO7JxtRGrXmERaHuK+kBbEiIJJOhhhanvrloicb6gnleL7P9JNGtwqhjjeVSN9yaOhzHypC3
9S/C/6HaPSRQ5a3xSoMYr6sW37jy40pkcywd7fS1Vi3aBmBArObDetyo0C0Dz4eLye6jWQKL6pU2
lHsddbpx3gAKJ6XTYWOyTRvpvipqWZx4pn5fEskhFIWvY1Rm3/Isx2WK0U68BH1V1WTCOAO8LKaS
4RkRoSnM4wvBNkEawZx1ir+NWvAC2dKzbkezXnj512VjSHwg2u0Ggf86KQTE8SGN+C+uipGPWNom
KUzLqoM/DaJE38ZBva/8fTxwSvLWuCA2A0Op/ftf/C+PuFWJuND5JAxBpvJq2M1JeqiNVpOPJNVI
Yd0eBKQhLdToDpIoip33dbbUhgrUirWgZkwXjvhHyey+rwISKablCcalu7TzyptFOMvEqGLF2dBT
G470FVOWIsc6nDRZkUFLxcTGO8FQPq+G/8q6Ys/C0iQNoTkTICPkcONripEiaqpt80FBRgGP+k30
/Aq4qALlOdYBIkOEpZmCIyoRrXn9B+GocbfwbiBQE65BHX+/NTVHfT1QyyiOjfBZydfRKHNu0rkz
vi9eTnkcK1BX7D3du6HH7UZi7Xv3ujouupLEvyvLKuCAclkvD/IBfbn/Ak9S0TuKcCI7Y7uMD/6S
vqAQXPNBNwucnIlinLi9/A03j4s6QLt/hjHbY05fQeaffwBQ1QvV12kRyG/jEMZf2cgMAGwPJ/63
xm8aFkMN7AW5eQbwWlSiyTq4Tt2KA7Kh/IWEruC2nneShJ7ELxEWHGqQI3KFHWRQD0vfb5m3pzI5
1bc6Db6iUIcJ/3AL/NVPVOO7vpYks7+1wC3MPs+SWLSlK4Z2W/fIUXvIXIW/KuoI7V8k/MnkV0cS
rQyAITZUqN3wmU8cj3ipa0hWemqKj156afbbAlmNomHiIdMdrrxIFTXNI4TsTPkM6nDhsjAWcOhT
22TIOV/D9C6KaW3qNyI1/lbDRiMnR8UfE1Hsy65EWjkRux6ah4RMAMEYKiZ2n1INbTxZnWgRww1/
s9d2ILjE368Gqi+qrHp0/UOTVDbNxB3bu8LQwgJ6s50U9wr7+GfNXwSOYXP93AUUZ24JJouZLJQB
Gj+T+Prt50qjr9Vb0N7vFJYMjvuN2Tnwme5vCJX2NLp5nogUM25A394Ow0yK/1AKdcRU0E2C/BXe
QXPDH/JFahm20fdjZNWhlkcbqgT4qCO9bt151nLSJK6RR48YXVEHiMuhoN5hQcVXXtXU56Ar68OW
kp3B5Y8D6RRPHrTo8V5KJm6DW5qyR5gKb5HC4qeNdKypk0+Wbp2KfcZYRP7B9xv2ubiiEZfHzw92
1bTP6Y8rEmrBJSmSS45TaP2zqwzzLMFJQriW+eGK+3AMGsiBdNOsb8YwDLIO6fv1dDRntfDHaZlq
79SYFF+T8uwA9uEmt/7MGtp8HKAXSfq7GXf1uDkWup4gepQokQcA/rEHvxjaY4Klai4gjugxlipF
5PAeTXi7v1OJefp7Kj0tulWzMFFhS9g0upPBvhuM8Npy+cJar8SkcYEpO4RA00o2MpQknaTHeNlo
+FFyUbNrlP6/ViRHDySCjp9oGD2n1j5wu+wf9wihdHQGoksiryCnBCEVnyc+mWXhMYs8lq4bIbkt
HpNmhwyVQZcyom/Q6v6GvBEHgUswFzkoM3jgPa5sNnri3hlnkqRY/PGA7uQ3SEqQqiVPO8WGukna
JRtOrSCFPwGalibi0+XmzloPVbal1hoBbrmdmLSQIP8+bZIr6dzcR0tbkhQdMVUQZFvm3jhB1GLa
zI3eXDaRMj6bJE2MZKHOKFXxeTFpFwotI+bUEUHukj91bvvHfXV963Bfd+HV3Gctn333UxkzLv29
N/1uRQ6saXuN2Cbk9lZxq3g5gbwxxiJfSc7lGjaLfZcvxUYnEqp/66Ki2c4DcygBR3FsVRgzqV3r
I38iNf1LhGqFMaImmpF8eEw3D5AJoIlb8F/JqGd5v6jQsqZBfWOyyDyxILG75S+5qs9ouUFARh4m
Uqykoaaiyfvqru5mZ+5ApE3Z+cTy4FN6b7KgRRkwnv2r36TyrzBgHR3UW8btocmhNlppVFMht4KJ
SYYvNFLVvLvEyO6e6gY124cgQb8LdZGDHUCAvt5TV6D5RmgCO7D9/bYah4KrkhAo939ilg40C17G
fsgodWoydeKNEatEjWJJGHiaqRNlV275PyabdgYAFhbJSwaqm/wWareklFh6I8s/+3BqZ+NTLxXn
Nka4aCyu3lybeVWv4U0EbzZjm0vxZYjzOEBHM3cg/onK7IpeoiEzWXUORyZ8sIQvuJM3iKFXuYfn
ElJ6lcpsdrrcTLEUB6KXy5/IdLz+Z5+wj5yCnHMju1peO8QbIfVAWTWouNQXn/+m/+awnK/RwLbj
hOANEXBGaYATerte3ua6jyASVy4tAQ75SV7CRlYoGtSidMGhd7Cw+6cx7uoGWp7CD4XfcynJIvxP
qNBrAv7VjHD4FvqND5qJ+L5LLwp3Oh0dZwWWYGArpFeejl+DpOV74ZiqmnpU4AwKsnaYaBfns/4i
6V9wFGWGfOT2f6Xji7Js/Ys2C1JaNr6n4MpGFw89e/Fv1ObsloE324xSOudDOcKv3TJT0klqe5zd
Axz/WxlnTkY4cSvJ6+m2DZsZUVu2a+xLzRJTIumPHsF+vwTdpBzUI4ZBsGNSRFIygKJoJKmUraS4
y/Iic0TcKnLS2QFTLbENnoYUbNYaIRtgVxomyyciiXiQUn/5e3oMVrsxsGaVFL59OOkrSWTSUiKh
r17sXcuNk1kUCTQ02z/cBr6bacydkDJ+ZhUOOxHPfuvSOsJS3XvOcAXu7NMF/X3/bwkaPm+nZaeG
eEVUp/lTqehqv0DLHnjnDAWGSMX5M+R8fU4E0nuwgmwegwZ3NDoCAVvV4kbujnJkPQ20m8D6x41b
fBB1riSEwfUiz5QZLVSlYPURc98f1gZFbfqokOXh2TOtS6wxxWk4QbZOwPYFnKhF8AoX/1ZS41YY
puuTA40AKb3U4lU5NK/obsKSU9BmNPB1N4qV+o+bbFX7IcybQUL8rsj/wYTT6Mql4e8CsWWh83Gk
37q4Egvh2BRookQlxN7jJkIyxOoE8odDUSoZjGBoy/wHcS1dF6ReLqyE0WULAPuu2TYLNbWIhP38
G63AGwr8jpazYCAO4KCuesMlnajqNCmZxeXWpNaNe5yjU6BAdWEL354Xw4kOYvUIelM2BR4mrwri
l9yp9jNecHWWCkCjq4FCLlD2E/wlkbdcC3KxfH8Q2RxVTrVGF86I80xKJibZLP5oAhEcCBEpAn0E
HigtjvhvAbKfnkJwPOJIHFyvRPEcJ+uFyM3FZCkl0DFNHqXc2bY07gPEfYAhqCf+CIOMbneBoCxh
u4n+FTasfBlCRewYTdJ9Q83kjvEr6mIreT3pe8Glx6Tqj6IgNuHuvVt4H+/ioIE1NUFiZQm7qlRP
WC6RB6G7JoFFChXVwyG81HM6TW+AMhp4ievETAw6hLFq6pswZ3T3L6OGZUZ68ORok09osfgkMaXd
8u3Qa2CpxQ41BJ4Jg0U79k2d8htUPkLbOQl4KZvVxIg9K/lYTfeCsI6S/2VMQuiiwt375g0EE2WH
W76kT+TIFZ2Y7Xo6C/jQLDgH3WJXAczg3vs5FOW8MkxViK58zuUO2Ub0/PCKc2i8QE6IAuF/wb0G
yqeiBEs+QSG96ow4SWBUvggSgUXQEJPUFbj5+YWts5J3qopiR62vcf+EiZOGdp3ClTV1lQjw7Bev
7i2g0F14yvW3fFI0MCwpVtJR6F/QprfU2He8bdCJH/yYQbs6io8eo2uRPcaBsY0VT3VKbCUdqWD8
VUyCY9e5ZY9gtQEGX0d3T8O4LwrCbs8BLa4dK/YGLz4TaOHMJm5CBh38YohW4CiVNyiVqpPMJ49x
O5fEcHku/G/LGOREQgBWCqNVvFGmC2aUUnl/vdJ3uJMiR3UYL3lHo9LiVstRigtTAMnxt4oI8wA3
jlx6NFDPfxXa0lpgnM3HkFL6ctRXmH/6ESc6yXvGn5oXDT6w14wYgTaWjF690BpFuMmx/+rz9hwO
fGDpEt+8Pzdnx11JgUpQLvobppRKpDrobKCQmv15x1Eily9fmX8QHcQjv3Y+KFJgqYWpcRB84wRI
1ruHyogtyIfybNCOfqLiXSiOw5az4eSA1G+qwnBJDXylLxhsYUMVSxuz0e4nzPemDczzveeVwx+A
1e0SrTLhvAvsropzBc7t3YZNGAJmmTKzNe52Bw6voVwtaWCdA+yMgMQs4uSOT7g9OIMJYahlPBBp
p+YHBfVK6yHO4NefnH9yKmS6r+zKLWq1xA2JhxqR52ZCeDHd7w7WtbtMKM5TSvxaKKXBSoZJ2b4O
KpbQBju1D1vQhNeKl659y1pIl2+drR4+S2TQ8UzbEmJCegdCx3k7nhm2DtXQF3KvO9Q93wtHuRZS
wzcMzKhpdpSGe4WcFr6Fwh3NbersdPKPt0IPhHXgltZe3YACeJ0ZDrhDjZ8Dr1D79dLw4LTNIJ6E
Vdj3WpbVf0q32rxOTsbcQaqdGwg+S1wLNwliKvKxrQB7+GcaFeKVC5Pc02bppK1p0NgVvdBptJUr
Uz3dFE891DHwBYTklEtN5GVgKxeGFd1oYMquN3d/1HKmpsrwY2rkHrq0TvDcadXEVMXzdatQws/T
XAGQxw3jGOW3efOLAaDEZK7cB6E5rj/uCKChTSxXjeq6LZz/7c8ltdyNIAfQc45yrI7123oBdIOh
gaGqfrU5kWgtLF0JjkGyx42x8FMu1BGfkaS75n6JJwdvkoIIp2Pwgb9RrgdJlVCAqjvSMt1zIiIo
VXMLNhhjB+5fnqiFlZvnDUcXwmTqQS8+paHiuGbJbxOtBOnzzMHnqbsVxo03QoWnQuL9JH6fPqfv
rL4o9+aFRw8b2httHCg0jm5MVsoSdTWdW1+xLNgLmbJJccMQVFCvTuwr3RMOvm6M+fZUqOt95uqF
LZi2TUdgyZseX3pLp2HYrPzJnAqGWgTgvbNJbYJkE+BMJGyWl1mrFo0YXttLfeyqoRwAxwmNe5GK
ifEwf4R2weLhLAPq05lEiUc5WlyPmclA6IQTHKf8AnxZbZXayYagSib0pnHBoBaQRoZvVwEKnvgD
of5DB/TWLZ0e2CdGGjGIsQ3azBMcOUQDmVyQjwIRVOsLhujDebBOy8Q09qwxoF5rSZ/LuLOkGRtB
S2Xlk6uWy+4FpSibhbJMOu+xJOP+cAa8dK1fZxVEpc0qA0HO61vU6LTPa6N/CbtvflIIOLn3WdKU
atDBWml46Hx11YaLeIrW+s1yFVtGIN5cgwNWbUZZFtTj3jMsPi/sBNZ4mEzS2UcZ2/IYJir00dD1
awmYrhbhvrfvxoYZrI715Z3ThHJZMireIGxsnsxriVbk0PNOQZxarRTGBMuHFIabIS3ADGBns923
XKM9sF04fZy/a8ZBrBgOafazoJb166THnsh1MSiMkh+CLeZQHHaT2a0Zy2tcwHv3WZZA5oJix1KZ
qkfJhmfECl7ife+O6qUULuAOLJ9pr3vSG3YdiR/vJUJDFPoPUbVkw1cqHTrK90oPkR+T2c9HY7kR
WfH8enpUa0ZRR7HWclStJu2ELxRXtqYVXPoCBoXgdla1nIYmZAp7DZGqfCXVXTqPKrczKnkslGG0
oaKlZzgibiljj+YvnnQvWzUqplepCBlSKj1g9vBTQGAW260oReeb/2OVrhM2+8ghsJzXkB3qosVQ
vO0NdEZK6Ln2RzRCELtklQfEu6oKIsrQQLBk5nue6UfmaRUvNNzEKSstEvRY7mAe3lnxKXMMJVtb
BiO1Z+Td4pWX/1rD5RZy9XGbR+MmDljtfa5kOJFGudvsHjF71qPQlP48rQMIzrYhPokwwT+V33ql
KjfJY4FicHpkhX5HopE3hQrSL32wZ8DqjKa0yzZYHf7wjAi/K3n6CxC5QawzqWN1xEX8622FyBWh
GlbaUbi/1I5DVBgd+B8hh+EwXoMl8s9cqe8YshalbuZ6uJLsvIN7HDWWNOURgr/Aibxj3+eqCiKa
DP4i2lmksgzcDkVzLWHy//2BHq2+fe8cUjjA30pTCcJltbhW2FlshRlcm7odEbSaBLMG0EVqr8wq
vF8sD7G9ZQJDV+QMpkzj/AdqPzddjkxabWwOF1HNIbscMJNloWQzGAwxalhqZ9AB/T9stqGDQRrv
FY0JVcFDkSB6iO1lpOwVJv8B49ViVD4zRODJ3e1OjEFvj5qzeaS+N14RTFqQn8KHhD/z87/V+V5h
nGv8CNDkQfEeuVPsbE06J4LaZUvjiMVFDsqrteuEyToM7vmQwoT7VhvbBppy8kw3yk9Eupa2b3PJ
bozN37TAJEV2k5H3uWkLR/LH3jXuG2juHPee3ApLJT4JyuVL9LVF7DYKFEDeJ3VXgADlVtyQcoG4
lJyJQPczbFJUU2dFqfk4yN9W0kX3PE9sK4Pd+42sNKrulKsUQs1mHZNM7kmqunVgat6nh41rIB3v
ssMYGowmCvlk1vvWRE84X2cXx/9MAywIvkhZLwziQx8NB+Hf1mgoBa1+LvtmXn+PssRuNlQxZJx3
ZKCfsk8PsPQFEOpy2OoASZcCQW7cYZTVQgmmzjGZr/O/8Enkvz8hlLY2Za7DUElgTZGNQHKO4Udg
S1mar6ujPt3tcykvbb4IyyxQXRF+8uEoJcEVst3e+cxtlkNcD7Qqhccu2j8zSPQRUyxJI2hWXFyd
cRLlfCItjQR6NMTmfoOU1u9DOoZfjDOPvPioVN4iQOZ3pEcQbjH+RIcAuRw+W5AEBWisTXxVT0Ve
RIKcVaumNjI9iHve6j/N2bpgF4lcHku1YKh3TSvbPc/rYnvGPMEUiqKYlu4AffagIySmP6IiwBNt
zK+B13VdL/up7qtjgY+Pl2pl7LcY+BDlH+YGbiFqxTUb+CGFa8p5Q+8ZxNBAsdR7IsAXSnpJPn9f
5D2wAUofGqmXriCMYJ7dEZ4uuxXvv4gltyCn2OMgUairWwgM9YRywA8zvw+QTr/TPza7/uYNzVI/
4Iti5LoqXk8U2bGCZO4X7M8dCt5Wvvv1brL3pDHF9DxXL0qkme5QaOhc7R3UMJwnGEYKjVuwK9cq
Q1BlxYGZtwQN95hbZrhwjH0C4moDXDqAQx3Ly715jlHVbvmy8Scmm7whQ8V8XWpdPuHomXGkziNO
a0zcSTEMO3RhRA+SlQYmq6gfKCkg0+aMaDAhEg5yU1p45/UJ3Q3yFFe9IA+2fiqw+SE3nxvyCVni
Oz9Rrr90xUaA+iQkqso2qtLQ/3+9LGYsI3EceunxiaqsLN3Yk1b5HW/qxS21CdAFJ+jz0nxqKxnj
88pFIHzSG7RyjSPbcB3zZkpoLQkq9t+rPbbkqwVgmbop1XpFy2XCMZijUSM2ZRQc5KscpzERxdvc
xv8oqvLtH4KGo4qYf1oLs38TVR5SvRXyhM57i0hs7R+ZeP5omv20f6zVb45k9zum7Qti3zv9PEQv
mpVI2usGDSBhWyOQJFvH7JmqbG0rLkm+W51cr6DHBsEIZke1EJ2rmovYXAnPcKdoP4ccvJ/W1iEb
n8rLCPVg+xSBK5g4cFFrGaw97Hr67rYpSqvzGB5lXNAUv/+TrAHCkiztEosw+lEnf4e/HswcBpjA
2+3D24iemCYvV04CbYDdLCKFRTuIEWePc9xqB3qJPuuou40fLQCO04/C1HJ3p3VU4mpcKVx2yuO8
ANIKOwfHrrbh6HcxN6UAdhMqu/PHikwgvnvMyJq7MVf4VOhVtclKMZQCtpGIBpZJOtHd4pHHmrYC
zIdRXuzreO29YN0NvTqoMLf0WWiqBdjU2abYhE72cUaza3cnVUxgvz4PofEtHq0LblDUf+JPyfAQ
nlwpUT6OmuhWOlWr4fNLFHq4NPo0HCIZXi6Eqfal7RFu9Sp1bCl9ho64vD7MNrr6+p9cpQlbZRwn
uMObmvx6kvCeVz5QeO4YmkHGXY3R1EuGu/eJK3FF4sgdp3HUE0dhtqUel72adozrh8H5jwtyld4i
EMfgTPyvsjs9bYoNrgj6aJ2ZYEV2GEXkPozZl0tBJwlHtIpVb/88E0L/Lljvkwa/0PkvLENyToMJ
hpYAAqu6HajrHbsnb1YCvlC99/korDMhivoU8TLpca+e5jqvxwb+i/0Pq04lzQmiJdCuk0qyRuvN
uhCCr8y4EexjFPtDdW/aIF/j+CCOCBXHp/c+53at/v/K58R11mHpJTtdAMrlCa+T+a0F+UTnGm1b
40Rie0m21YSNx64N/tdehbccJh9IZa/1hTe7s50seKdUSmr4EDFXuh0Knuy6qAI4GyUv2drMszAk
0w+sCW87LaAox5NF7rqjfXZWfvk5FBW3H6iqW3BOeHV6Ks0JOvYPIOHbKLL0ShV5ueSo2k01fqkb
B+7KKHZDZzEzz63OcFrSIMj5+/MkByUCgaqby4VAbXLoB827X/bwYizK/nNWUS/PFTYX5vX1BiYo
mcxQwwkn3USEeOBjjPyZg3kaxhgBl5Ws7wh4AXqkqAHl3tfytv+12wDvYt6Yk5AseqxKEAgKx3J0
lxxxsKYElcoDtgttEyNtA3EMo/fAFfGXFN9VjBuUcYwNQOgUI6UtxqtG9udavsfivLWvEXjCWmsj
PeeIAuFWpEFUutEC29jEX3etIKnVMPr2TLyQ4Jn6mA3m5OHGyMeUOrMyxS0TYJ7/pLNWX8ZWPvRQ
gmtaSJ2qyUhRyNwsU3ESkmyY/m0g6NoiJrGO+4VbdXTP0Gzirkazr3xc7PFdAVeRnq5kyZJ3YnvA
AKClUhfzbvgrlCycdqiXUNhaIo1E3Gqo54YGuIsHt1oVEf+rwgOsXJiDE9QEWcAWaF5dHIMkcz1V
368i7lx0+QhTQmaXXMQ9qoL5fS1J+G31u4ezQc31eX18j+LOppfjGoA3x9kzv8cTJRAyVBlxNrFP
AicVTjaEMEmjaVurlFSUdp+AJez87PjSFa72NtteqtO21UDE670A/uMA2L7ECs1wlVvO0pNPX2ME
Oh/pZug9DJaWtI1nf3rhaaeQSZfoVjQ78aCL/DfRNCHowBhlv2qTWTDzIv5fgj4yHB8AsUm4PC/Z
Aw9pGw0t545eFJe+08NcjzexnP6M+zhohwRRviV0+79Hx8UFvhTZw0yKSXlzBYqXg0L/zQpOucV6
QNqPZyT3POaAef/Hyei7Py2vvbC12ccgEcRQzRj7l6oIDndnSyq+fsyY6OP7B+D1HRCJdt/2ot3S
Pwm4l08XvjThsYQCz8+C/rY+mlPcjqtItkDY2LP0tQnLIGDAB2vHnYsG8i3RAFFM43bhtgAvQUzs
TimEXQIY1OOywRtl2cNkvskGMvsFlkWBxp5RC5SFzIrbl8NoyCzUt2NkomqWzBFjw/QxBFZJhKht
ZOZkSzcgifhAqOZGZrQ/RV/XVciQqFQHV+ANKmk71Kk78L/fRpkaTpzyD9p6zGF1SpVzSaQNXXx/
PKxOCZkhZVueop+xFQhaysUMfZA5CtZES1ukq8xVWQAkKa2YUYG1TRE1nxWTE6Rsygs6LTq+qHSu
SBgZzFBVxwZHlBR4FpUeDndA1WrTBIsUWW7JhHYl1eQLnd59lfSAXHfgcRy9B3uL79W5VVf071Qs
XFruSW+DHmQsi5bFQJH1Pk51+Z/Sjj4mNODLMnhmWdKse4q6eLOdwPJtRLUpCM/oGZjbj0NHReBL
iQs/a7zHOSWag8U37xfkavrD5pDUEibawnb6GJVa5Ha5kgJgtIJtHaq/37WO59W7dw2KzK0Zklc4
tCIpYG6XF2IaZ1zVvK7ypLR0/y/Jw2xEd0KuXG8TvEeynq0zcYazXqvyiLTX8jXzHJRw0Iln1x/x
mu0xAYk71dcD7t9ZxT5qff6sPUIScvpNU6jie6RRLE9hHFUgf9YNfX7rKwPajQKKMwMNuFQVu1+e
ab7vSkoyw2/B8iO0SOUVKzpHol9PtObTQxejDQ/NtLdPxpxNynXEawLa8p8IkmssCLOMyl00Twdf
/nnyizxYGOdDXKJO9qfpQHM2HTJMa6y6M+MwmXjkfl+/lHn4VfCBBkKMnq9Hzizjmjy72yuUchlt
tLqf3S2hfRPpWWTCnPSzVo55H9mfLeimUC+yn6LEkns3qkj3OY/tBUx0k4jDrTSVnc4UJHMtkL+a
/13FN9aqXDLKTTWubWKvWKK9JHg0LcKPRGnZiubzphsVIaW7tccBnWNC/x8s9RcdNzgCyrECtZjH
0GdpSY4Ez13xbS5ht0gX9dDMdkSTzxM+taOHMjHW8IpRXWVH1xUdzJ874WW3nSbCWiBtSPinpM0l
ESsWXXmPchr53NDR+7XdTUTNQy1lklHefKZSiV5sBvGDxyJO4JxkSrT8RtvsgK9vpiKsZy9IhGta
WWOOVygbJrcenRvvdieSL6a4kF1hVbOgiU10WsZhrVuk0Ti9k9gikyU7t77En0/E0NcIGxFvBQRz
95z+JmMx1ZvfOBU/EHK1deqqChkUHQnPS71GPv8FEGv6bLTo6P0sMsAJmOEm1mI9M0wWatw2XMa9
m6VtaA5CajxYhz3axyeVOsoygYHqjRGpT8eiM3S9nooUQ6HxJZlIB8r9VqnspNGIHHDy56T/4wa3
zL2cFK539OqVgmfQAdWLXsigKGAYjCRZ7KU9j9L0JZQvYFK4jEU4nRipTRBd+if+IUoikndl1HoR
IE+uUmDFkT5hExnqGSmz/LsnSC64a/MnIGE7ZxQIt1dDT4U1ct/6GD0NZif0YI9Dsx5xjhK4R6x6
XNOJzim7R2IBWQUjK6U6OQFIiP0K4g8MyATJ1s5GiCFGQXzjHwYZhNRH2BCCg6UvYEdwRi1bXpgE
ikB6sduzViX3L90bIaE/rgDuHUHMFIXeeqDn63FpqlU/zJRapgb5tUQTB8+rwqn419dKlHHMxvQ0
BQ7gniJe653GeXqK7rsprXokm602/QFhdRePoTo4nMwlDdG5ZmcY6uTfZk9kNs8VjWhwUQ2zzYas
/e0XYmG0k8H2SXNKqC17pq4tlOH2mrtyaVu4WaG1eNMn0jH1EC9KWsCg9gBUrSTLJNOWnQ55OW4k
bQjKA5zd2xRWfmTbYbUvWPqMvHiw4lmFGOeU9mjgrfKQuj3OWV2uN4hIX3Co57g1Axg+5l19LXIg
OumHdpSB0MtsLIwyQg5BUc95jZ3cjlFhqpfFpmW3YoJbjWlOyDTrXqwmIfgczMgset1QQb2UC7t1
xELg5/xWPjm8ll8GhH7j1SodVU7oUynvSqxlsCFmyphZIMlSZzb3ivusGLiV1PAM5d08MBp+Wear
022LC8BPZGmimjkmZ2MAVktJ4VVAP3rL6M8KasU9W5Mzt57uq2aXTgBmaqsznQEW5EbIGTIn9vgk
Ma+IH576VsZdKWa8EC38BlgkKDPnuIFmRltlCOS2h+szoTlIN3/TaEwBjy32ffq+tQzGHcUpPVXp
AoueBj4YwvdO2IwWBzHiY3eTTzVlOA116+cTJLBXxJ/BKNAWbktBMzMnBWZ9RXqrkHmVdk+lkza2
ynfWgnZhRZgaKVB3W1jslUnd3SmsdruY8NZWSC/as3enyhQVpgiBqSYqxlrFzu+34AUVdaavNU1j
O3Egmj3MMc9UNGysfs21pjU4UE54kBGONWUYCxip2WV9dn9KnFjrbvzqGKUNkfnv20EHCKTEh+FO
SaY2DX3gwUDiTTcgXJJX1sa9TTVdj7ewvr4qFQy3bEdUWPRkfHthi007y8RYxAe9IJu5ADGbsnrk
fnjRWWHCtPC2WQ7jARyw8GkyNLv5aa/gVRqvTtbMlSHMwEWTWUIVktX8DIsRIUe+qRS3RCDoQZ4z
mH9gsXDd1wmU6HWZT4M22fxIBL8ByEmTTwWHTw3pRLCO/xySrBWw7Kpff6Acy6LwvDrPm5++BqY0
YJnwdEHfT1GehBdymQw/IXkiJPBMcDyn89lJPLlZS0B0MOenv3BOpOvn66yrCssDt7mzqLCxwH+5
VsHINU3H4LOdhdplF9zX5gHrpjTiECvbFVQ80VrrdbnciD6Tc9c/xrpuYNa4hSETDhTiSUai+pzd
gPITsLZfA4t1UbihB7XJtarz2niLmYoTJG9rYvkNBtcvtSjfy4v1WhrpSN4G5GFeUkPnfPYmWVKH
3MeRADFMKhPw2Dg0ILq0Z7EFCv9i/oICt/1SD+M8ku7oeuz9alwlya2/tYTLm5PtEVN9i5MMO0M4
wbhgHbpyzmBTNZ/l10MyEPwfIW6c+Lq+KtthuQFTrXw43fg9bKEkzyXXTDQDOC47SuY15UtMcsSW
J11jN/+Mp1+IDmkXwFWYSTOVNKf1iOW48mW9OrtJ4VZkNLMKx2m5YAIAIFnPHm4xQugPUCGlw6x9
o4un81Rp9qVMDjYYEQnlKyrRLqbRFFRdtVSE5ba4xgkFZkTLnkEKMqZfOWlvijVCbJPy8QZkrDHK
LRuogEzLFS+YioHi3yfRotJL4SnrSrBS0bSJq3qKawRUBZhoNpCpB6ECTSvdboD3nfLoPon6Cqmr
Gj0Yef6ldpzd+6hqf6rrZDcqKN3h46iWEl8dicTMTHkISUSMk0iRj8/d9/nxfC5zeH6o0+ktNYmu
1E49kdn0MyrSAP1/L8uDIn2iFrxWKu1n2X5Z4kb6g/E6O973ThHZHJCR/uaWaDoBnXHJCQ6R+xPw
5SYxwaILiWC0vAl/5OR/kvmcg/DuNOm7IIp7hJInGl36whzo0PFXqeHUHh/UA/cTokUirBHT88D1
qeB3wwgXaHuP2/N8RXBHumOx0oSIVEn3Ykd3Xzh/vVJ5HdAiGVmPRKdPErEcMdwJ8QCEsbylgYRx
jY4j8eno/3aFDh+9YffCBZkHIGIp1Ak+bBYR/FJos0UDspFjKYARg1ieXm5JspDUi0lc7zrVlCPq
EunGXIcYH+67lWFvZ6aXoYUjPKK+Pam8QLLsLTL9OYbiWDFIFIezRV4FTuenaMgi7ML0PEZJJ1/B
RGBBPRzOJH98ASFcpJVi8zoIzrDDrSNge88Mo6IvJuTV7FOjgkvYL+198HO4RDgTai7VEzbYEMwm
VO7mtMRPn4myLnLMJDLD6/IZHs2nR1b6ekMLOc9ny+rCIhvcstSlij8uYM/jKKDk9HW0MHOQ/Vzd
kR6xMsKGSGIGxAmMZPmK+jKTO7SLu5w09VcJDgsZpV86wj8qpx1KE2sIDG7A+ONo/4YwDp26Ms9v
ytJl3eVYexBYNtwkPkS4wKOCsnqOi5Zog0KW/NKIsXKgPWjJ6oZyU+jAanrypxPk1NVtdn94n5uv
z9p4xDbe+SyEX2gFMRMkJ3AR27sgcPvr5SxXmIulG/hTOfD/5qs311dMK5uU2VuzoNmVStNAWfpR
M3rOWeHQezkC3bUguH8yasbE9HVFNO2ZTTWtlcN5z3m7h5+iyWGGIIzAPNtPo4LITa1r8WZJZit+
S3/I9iM4rL7OBZZDhmgkxokOoRL3+c4+Ly6WklNgMBSFweDcNAOjzi/nlnK5uH00bij78UGPf758
ao+R1MLT0p76QwvIsW1qLcDLjohSJX9S3BKY2GgGEjjuJgP3xF/28OzzIhMzv9Y+TpGZpfgiXIWS
I8xCGwDRl/XkZsI1gDOa4gcs8S4hmI9Aw9RpqXi+XrHv1co1CTvZNfcNv8exK/KDFB2ynvjERG9G
pmTs+PX3CVFXXLXrRVnQUi4ZbbrcxD8MjSoH2qAQRu+HaVbfMvITj630+BHBBll1Sb+TfmXVInho
3/vuS0Ysxz6Cvm5GHr06K3JfBQEF7YGsfQ2W5HjVX6gH+VY/GgUtSL4rnWlmxlpQBvl5oydckmkn
DnRbtSKJZ7u4oGpcXQ3xovRXwhft1adH2ob6hH3qHMb+PE3dRcg9T4rkts3AAkmduFGK3Sp/GbAj
UG6C5zB2W276BMLbmZh5N4JsFb1hTs5aiDHCNvVuY/kRQ56Ef6MFG4HMEyK9gHuGKsaSV42jDScp
YLGyEo1bjljYFp89jWqcCTDvPCp7HUm8JTnHLY+k/MXTmYFcEAKHBzNLFwqYN1/W+Y7E82Ebrfro
M/DKOHxjCk8TIEnFTR0YI0FT5imI5H6cHB9qiy5UNy0I/FmARBqCGPkdEeH3ZCXFI1tnBQRd8Qm/
OmO3jnDlFNjeBPW+xh1x2l6PZ+72Y/LQ8n9qvACJaWfQddiMxo/9+M5wp0Tc83UZjBALT+C6eID0
ELx9FbiVLqJeRzM+EAzGO2b4mW+6JrpfIak0JtBWOcAcd4ftE1kAxUXqI8OpypmTc2o5QyGsSp9W
SbsXDfAXCMIOcyfmrjQ1RaE8ZU4OmWwuSXnyZKbA9ULhPL26gL4cvLDA5yqXHgV1nbkHOrKiQke0
OlI7ajY63yTAWMCpZlmPOSjhFbgmMnyQQkmByZvYVAM02pBdONbm8UnosZQXRPDHqy3wS7EW70bN
yzmiMTmCDO3ij+9LG/y6F0cGFHLa8rEcO0o8O0FsCcfkZOhWUEEgDYdDh984DjQWjW4SkT5SeTIk
vJw5Bzp79Nc9DJom+DBV7EZWwIPc/o2gjY4LaEnddbAIGgoDbqcI7uUq9j67sdJpMWnSYbEQS0YE
/yGL6gm0TeBBimY2Koh+7V4goWMyE5TycbZCKKwUIxWNk4D5IowBziukXk5sETbPhxZoA+jKq9xi
wYz4fZISMYr3bEr6TqQKe1eFvD+TNw+iAGxTH025kbXpPimHDjot7b3Zj09VWE+8K2F4ELOsrTE7
aWaEgDjCacH/VEmZKK7TCgHsOgLHMuHnkmU+MJB6G7XbaULbp9A3A+32w+BxQAhlFN4JRFx20ne7
y7zC2EseF/ulLqRqSBsyNtmKsJhvCfmN9p3CL79ggfRrh23D/b559/6T0Jpuk6yaT3Tui+5c1f9N
DbcSqiqw5uM+y+Dt9I5tA83QHRvKpF14lhRMvu4+Bhyp9pBqoEGD4X3zVFhFrYe4WIfH2YdYaKGF
A7WI+sQTZf6lsA6Za8YWCpBZXfjMAoK1ZA6gAFGC61K9L3Jt7QfIiNrvqYk5halBrwloSr/yX+aZ
SHur2/EVDffoLD2P9HP3Vt7SSCpVsYTekETO5TefIkhctkvRAlZiyg0YAJNSujlToaQRbWhAwEks
Pp63IXm2ABQEBEYHJBnmLteKwUssXfFU+pLSk2DqssBl+llwucu+2SNWMkCpJOl6ggcTI9qpGMkf
1C8X895V28bHhIncuCi6IwprTFXb6kR/WXVFcIttlavA1G2k8vZK7zV4u67pQXOd1SUBaKE3AYCf
WFIerMHXtFyxsAu3gcTdL7Mu1Kuid38nL8xZJcDCMc5DHOv7sHwXMAh4A+podJppVVZhAU/reUg6
Gsk98x97F+hsZ7Yww3PS5XdmXAwZdV2Wy5qKhfzAM+P3Xa4oN7TXmu00rr5VYfPU190rERhkS3qg
v9lbnQ16MI0g8BQ7oQDDQvtiEAPdKcpRM9cQ77Uei2X4f4E3FFe9m6AJqiSxYVdrHJQd/zDHPAfv
inmbwbDSdFVMSa5w+HydGX5NumgjWGrGB3sAPOOETIEnZby8ihg2nQ+OqBUJbGAMTTXjR2RqAKWh
t6IpnZkTpAgtKd6K++1sIm9KNncvwb8RviB6HJ9hkD0RxP0Dm5wdrwZTEaoAqnVKk7rGsGHCPfPX
6sjF9lkclunEOkm2KFC14IJHY45Wucoht0WDIXzGkLAsSOOuKiQOL66KbmH/6HshaHoKkjnoUEcS
MrXbcJfuPskQz/lTKb0Gz8MtfVPoGMn5Lq5HCQw0is7H6BD1OoC1ogRQT54fTZCHkC9OpomJYrd0
h/WPQJ8geeKI84QT+sKtMoCabpqo0VoJZx1HAwTsSAWTI3ES2ZSHjXK7sMGl3UjvuNqJ3mrsUhhN
ycFvFTdCUWCmhxUkh0y3miglLViNNzLdHjjKBECXm6WPuRWsoFYZZXM3fVz5QphsHcWBpmtjGC7Z
DxBNGcNhRpgVKRFfFA8kRWdkC0bmvv831kiEQSU9s2vuxc4Iv7Dir8jjQ2HbULwE8Pza5mgwM08p
0Lr/jUqXsRW0h+cTLoZR3Ctt/GRJfB9mppFsN7DW5v7QVB/LfiQ9EI8pUNfkiB3BFbFKqJM0Tuz6
+x6ArM+b/IAHLvCyWojGvXSv3qvr/Hbg89YSqvtPLfivm3qokiPl+gGGWxQKPZl/QP/B4vqu0jQm
qFHhAwu1jlGbTNGqWHFVJw/pav7TDioGsPUnWw/sJ73e/xvGbiC+SppcekId+txQbyWcCP/CVPQR
LxZk6H1j+XT7M9je7v1TRD9/AiqTnhr0zZBgp9EakNgQ6XSs63NYO8SQnIHcUle4FR29z0nKTZP2
c7SgGdj+w5ws/ffkT1VFQBWkLIx4Agn6BnDAqHKxipk7Qgxqvg+KMv48z1OMk4gh2r7qa2MzCSZ9
J94sRlV8ifB3H+/1HjCpabnLNzNheTtMwMvr5ue1Sann1Oiuc5Kvfm+lMHAH3kMB7vayKO/YwzgA
MKl7tEd0FTF12GuiHjlYod/w0jw5mpWuOYPZGESLJCp/eqVXWvVA/HVLVd4kklCVDEAwDjmz41//
MicWhvxTMz3/+lItk4MrcQvstIV8FsP6YI/kw/rklgvJNyLhAIS7djANxhzqHnildbnSu10r0gJ4
ZFvugPquEgg0Tnj/bYwkdw5nvGoHS0vsXQouv6yp0yzfpYGA97IkZ3WyJTapofLk6Ru9kRUeN1qq
viABgUfkcPz1BeXHueEfTeH8gA28lJZuviF7YKaRc5oycCwChWrzSM1mlP3lsyw1xzaSNxOqt9wd
VCgg5AkLelvu7o0JB0bUfbnitUCHnYHKWWpB9TMVECDWyBS4wV8HcNOa8CbQ96VqDKAHm82VFUAY
WCyK9/nrymf6OWWCdOrxbNe0bvZfhhghmrfVZ9mj8RFdObOavwpx8RnlmBT8t472+GLJc7QT/WFo
N3OdE/qit6Zf4O8tA7vLUoAyXzvWOnyn9XirGshbVd6QCzjXzq/m2sfQR4modROQQ6ht/BLBDuSA
aehLjf7G88DBdKDg4CJk4uxq+lvvb+O8JxQm/KefU7b/dbIP8JYnRfY9jTcNS9LQTqIbhFtua+gO
w7OtQdhq5kxE16sp8AiUeUqIOm8b5GjZryoYUH/Mmk1moje3VcBe3H9IVq3u3q4OJ3bOtMiAheOM
CmvfUCY9OVaMIhJGjrUrPTDanjJVZjKetrOAS8oCGq0nniRwvO4OoFmJRaA1fn5LuSIUs73K5PhA
cSGVIcANfJ4kUtNkirnag8yzrv6TzJLkFBA2fqeER2m9JUQ2bLnUgBAYYsFpgUGkcVm9n2626i87
h9lS4J7QDhQrZHBy2cYgp3ERrwGvbPzpLfOCzBCoRn9gF39Jo/kWj9563xLdh3l2NkhlFYdy/jc3
Y3j/qBM9D6i+aSnYnDHlMykIRo1dzLVhTnkOc7KNRokZb7ilZe8HxmkMIfBbUCP/GngoyF0R0Q9m
lFWeGZGzma2eJOAgpU3WANMneZp2BauTC/mOHc6BNb316FtwM3GEaIPKM201knsRbyTmpjNFBM1r
obhqvBe+mjtpCXjqWjMEUal9mwFigj8C7f6uX8kVy54sw/F31/8pikd7PNyjBiqFr/yzf0MP8ILG
0QjL351TNx1qR8nOHPhfkDRC3nP1VoKBFTXjxZjzSnCk+r109rTy6qZmH41hdF5HIUFlndBEFqAz
YGRPskG+wou7E9IwRi9vi75Od1Nj422LEWh/WXS+9bzD0CvuxIfRZ9YVaVzby+riS+vIuDpmPfXp
ZNbnzWEaSROCplOcjaN6YPttSGZiaZXF0CBckaAhr+VT1zeAKxdNwJ1T73t7Rn9D2PU1CSaUVI3l
wZP5Zw+FSoCwzYnhXycRb9DwhC+j+D9jit1T2ORwG+D7glul1loldmjZfeL5fpdgh/7tULguwlgS
BYqudLQcg8e3FgZmjIgx3+eTA83C/LeO5L+KkuvWTN/sOQD1bXOcYBZ/rZ+60F9A/dJxCTINcouC
QKUzG8kEZz1vaayaAH90g3Q4XnstQ/oj3oYTpq3RSfHCL862wr/1wZcC+KBeaoAUyNKKjhSqfts2
LTBu1OX7NVPXI1X5G/js0fM1N9bZmdM0RcjFoOWmXaox5wRun6eYxp/iLxPnVR+prqgdvsNvHYkM
D3hwr9cayDAWl62iW8CxBSd+BtF8/P6DD+Gj8UaxGLr6tNkFdYquNj3eePapXpEKFqlk/Z+1j7Rk
wZG+u/+r0+e2OVUCveDg7a7OMbWy/jBH0yg+yuBnnScCyLrnsUVueWEjpMMMWI2iAkPznn/mSoZ6
vH4z+v/H3XulrlCZLn2wchoAQmBzVtikAU6+hRFkBGnyQ2wu72jirdIWhTnMnRcMajj6Xtx07Y/M
c8q8RLJMxkInc23NP58otEfgT3RQbWqB8PsIWwL5xLLWoFglgo/ExcwVb2wGE4OIFDQioJALZmjG
umQrzfFbDeV/mR/mzPo35iZGm7j1H/D6KcwiqxlKzWf/q1xnP+acud+YxIyDZwC+WLzDxj/MNy27
vPl0ZwvaB8imc7pT8uJmwl7xzP1cToQ8692xsBQNkSenYw60zSd7t22W/OnCoZxibvSCJ13fYsyu
j8HB1eYQbyClYxOomI4E6NktECLAHA8wBpbtPt/YwBD3Gd9inwFZjAYByE/Id8xGUDnsOImLtQwh
5efORoolQAA8/wablQbpy220Fu5xlCQ4jtf5BTxm0sag3AVetBSf8+DS24uKtj7onpYR6X9vUzLW
vybXNaK8UXuBEnd4amPJcpWI10I1b6tZTTwKukRbcPePc2nfo5cLpQOpW3ENBOVp5zScIO39sZBH
UErruZQdu6eJVbqOMtB7PcuyYCmiBjvcerqTbNo2Tw1PiTDFJlj4QnzHTZYMHre2J78eptQDUnMg
kSgE6F/UEI+1FOK3xOrAXejpS7eZjPbkdW0pPGBXol58OGRqfnFeBrjpz6/dN/a5DLgyZdK6zMEJ
m0vXwx37Ipbdp5G+w17ZToGdZPwyu74aPbWfrWLWLgjpQzm/pkj3j3jgichPWpk2C6K6jcdCCmN5
JrCOj7hmy3lYZ+77VEXzesFl3AhV4nHYi/tQrUmBChZAooILquLupfcWQrrsV64GJpfzCxXicqyq
oEkLGyrCVC8ghLp03cENUSr3y5yjSo2pk+Bv9+DO/UKPgtY56XZ7Fvs6yG/+nNKDfRWLPL/+5nMI
rMuCP2fT1OYZLnmkbXdJUfKgYxKsiSqY3XCC4HI6fRczqYQInm9y17LyulczVZ1M/LLH/QkfrXe3
KkBq9Jw3lH+Eh93aBz3DzpMUvACxC7mClWBIQzmo8TUQufR4rf5N3CJw9A4or48V8NeH+MkVf1QP
ceGlh4Unl5ug5y43OTPfTO41aWpbPvae/T2IzsSRBd2tvhn7K+dVw1GToGgrjstNeUTnNuBhbGYY
ST3in0zahgkXwTRDE78Lb5ZorfyYILh8JYLMwafgLzpqGvIoH6wKArquJcy5NvF6gSPh1sKNN8V9
3mjtl9jMcaWY6XJedPCcWJbXZpBA0vtw7xoS2ns7mPUIwZ7EAlEAHzN6daFccxg38lkTkKdSuyo0
oC53DUWwJ1YFLh3eN3GAYdWT2FW4N9fWLNNILz+Cx381PD8l7sGc65oZfe8moKD0IHz8VZEjT9de
Z9M8og9tomY0XWrPlC5NoTZY0zexDggL+nbfwRK8WDZTvoddNjY2S2AMo4aNNujqrXy3Pj3s3NTO
X6qTQ5n1Qz/QrQvkg78g/HjF9epLmsHPowzzAGy3uSizRfGgThlEI8izBloSc+Le63801ntWh/j2
lTwMkkzVd0IC3H7G+gIgMOJDUUpMIy+ykixGYpk9H+6fwzMFR7L/Hk7ISaBvYwUIUu3+2rNQOUmF
gvL0AkWtRj56Jcx++DXO6edI6K2ysgZaHlK/aGGFDdOji8LmkdalhcfmTGhPkViKUeJoW7yQFpLi
tGUZT8eCtf7NuQMX+L2u2+M9Gtf9fm8r8CwhJVEY55zT7GjwcINgKrHEUiL66scPJLQeZ+b0HenT
s0qrYfOyU30Ph3zNtK1ZU62N5y6zYMeo5XbbeFSQ7i7c8m5/2UJgY8t4RAwBVyJZcx/sSSX6L4IK
wyVcDCYO6mnUARTjbBFOKDt/1J92M6hon7UoVTgs55cbErbpGgMPB5EG9klH/vr/Unj9v3FiKdRj
v4c53JEro1SQDNR9GpwwOoJprxMrhxtC1ZYU2rfORgGYIBmrDKV+06DbfGVD3us4GW0+KdMR1sDl
aofUoqdrd1Nl5Suoxr4M3NthrIxPtWAEKDDre4GxE6W7+jp9zC3mZzMo6KmeboehFyw9GwgjiHoc
5v0LI8UNogt+VOmPtzJbAjbbtZIBlKknPwAyzV/cSLVYzBlF4igmDLr6k6byMQglsK3Vyq5WQot5
q4bb9kuXh1RNbd+SQPNYJalEkwn4MgjEF5hOF39JaCMI2TydqtnzNpqzD4ZvEjlE210Lcl9UgYKQ
Emvhr+4QqmIHIzb580tj0M+0gGyxh6aWDbgLrUiNNnc8WpBg9iyRqskT3QQw5UkvE33Z5shOiidm
6HfwDvzuknMbE8mKdlOBVqDgzYvzH06cpAKp2V+Mx1ujY/HBmYkegqCEWrq9B4dQvdFHYviUh+tc
SUZ9NBv2WtMQbnI+c5i5i5jS6pbXzlEpbwY/3+cKwNG4Jg6dzxi3QmgXQjWUeNORv78U8Qkq0Vlm
qmJl6S5UDYdBU5FRw8yeGeu2/wysLdOMHqbPy+Kw3jazL0axdylLmnyu2MkP9rIKBQPVv2XbeMRQ
yrQwoJjg53YSidjVegKAdgZ8N/8N/P1F5TTe9XRQEuOcFt+XTgWaer8eKnCx5GiwNz03PjIBtAUN
zDpSvWW/EvF6p10gYjqqb6W8qAcadmARhTebgLuJ6+eViNbI23bCRMNCrJhCTOd6LZGE4hza2H8o
oFFG4kUgeDg1qocKaTBwCRE5CnJNrmSAN/gvagMl6TmnXSQSQVnb6CZ+2q8fJJDxymb3i5jxCz6H
3OBcOIsNLrCozhoXHildUeiWOcPqAsd+eUFRmTe6GYOblJ6n9euYS3Q6puTgzXtDT0svCZv6OHth
23kPSasLBZZG9wVNy3iWjqw+yjHcs0P0iaOn8djHfdSvUOUnwNlpKoX1ej8y/pennzdWiRxmtFFS
xQNUA/RcpsMwhFygjOfYepnsDGXNErLS6qwCquGRDnwkCPGujIDIKixc1lgEC2bjz3OM9NLnooZ9
IjGWmx4B7ZyKwmgDQv0iyVIldLxhbxyV6rha8kKd7EiHKATqJt8O52C//Pon/o6e7N33JevpyjfM
NBjJD1YUgkbVPOFJP1nuWnYMszw3aU9ImBLMI0ED/WUMp5lVIW5yxOcOZBnNdxURL5G+XT78qk/9
lPpy7UHDlhy3r9ocQdRyot3pKtsxdCNQyqPhyxXuiKR35zXmNZ5LGXxYURHuV1CR9t0lCQDWEKAo
6Gx1M83HJ3U6b18GK01OrgkGKmINZo64lYCSHfJLSjeLmd3/YerUATg5MVxBIBQZzfo45RN4ZLUX
R/7ti8uOBgnRV8tPhIZ1rxwGzykSOE1H+jAlydn7Q9cYBsysg29hEsnyehrXuKUdW5uaFOFLcRIE
AEmLffvYNktwSVAC4bDJBzKW7wioTqltu07UpxUqRrc2bnElJKwKRxGtKLXuCH1TdeCXBrymu+HQ
lqpM9nW+FmdGaedJi9JVHvRv1RUO7drYOrAtF4q+v3TV1Vj05ZmsrRP1hPZn1FCDj+nLbvnpoKra
vmhNFzOaRgKkLot5sjC7YTYaHsjDpjzH19B+d7ijkStir9wuKBX9kMhLmikNTxf1pFNQJTvYw1uw
EXbm98OQLDT9XyEiKlhk/sb4Z9FjQBJWO9l1wSEFOgmnJL8Ro/NoEHBLrvRHLaKVCwpckNsORxv9
lRhfFbM014Ww1hdaiyKSiG9ylKkNFhhQqCcrChgIUyGlqM0HrmYEb5fgueKBUbbqDQ3Lez7NGj9V
vqohzFNZavFn4SXVtD1fzJyXIwbege3CBH495rt3g7188xuAMYCL9+J+5oyojYkp7IH32woEUhnq
eU+Fk9VcaCFCsXZHpeN5O9V7tlLiOnmgGt78kuXT3NCLXa1wBkho/FW0emwm5eeZAFDeGU2x3/mt
xZFPtJHfHrH0FG4scEQFC0iWrjwndeQj3+9QmOqIs3gAhV0EfaDzsYWySZW9osswTiqiuW3NGNiP
KqOjIB0vXjIYNPkPAy0+dZNgZCthsmvZvVkYXttj0bRzHJdzw2Df0A0Vv4PYWoemKeZybTrksECF
LnDwyD5l/B7ncG0OHJxYLUjHfPzfnKsly0IF88aJQTU9GHFWBEZtDIogIpW2maUlzx5qw94IP37o
9kBOUzHKCPt/69Ow3T2Ijz3JaV7jHWdd+JJeqlgnEJi9URCHOGAZlVaA0ScHjslM5hIkiX0SvBDl
prs637WbCU3n2V0Pp5IKw8blFptnatNEvoRUHPR67WsNJ9xFD3gR5IWqSoN/UQEy65MeaaHOHCTz
03ajLlrXzly1ML1bbEm7laTGxbgDPy7fPGJPDISxrWkhouq1FDpo9Uv/7Ye34j45btMF748In7Or
APcREgqZcpXsF3hnKj9ffDjk8tmViza2C33159CQxIQAws4N93/u/NvxQ9Jhv3HtM05krxPJoJe3
5eeZIAZ7RfYdMdugMa8IoTfUx7DmZiLOYQSfIUTJ2mbXAGVVDbQE6xuL/jron9PNwWky2Yb9dx3p
F/AYH5sph3IBttQI3XnvNjDI5qoKVSdf8tOG/n4lkjsF/1LhLp/ezS4mtyAuZcqaE2JFaJC61gBn
cKDRFTZlwMVnmXrAIULic/In1oLKPxXZmu+oUciz9VaTeD2nX04X1KuNJ84l4zzpN7I5sUyuvNoy
Nik0A8IEQxPW9SRXHqlWlDIthRCOsDoWsNCUjFawcDgGrTPl4Rvr9ZXStx7UIx+pULVdRGjBnpTF
969OiY3XhY7pV8KAHGcKTJfx0r73Wf2aVAhCmrGDH4o6Qg4lbtYcZeoJTDP74PiXPYJ/UkaBdLm8
eIJzlSDnHW8xHg75nvVhfCtDXvTX+rFM8V5NNGOgkbzlIDVM3ZvrSSPGPfTFiftRnMv82z+keSWd
SCpO3ThAKQZnr9Lqxsug76JuI09ux5syi/NXJSub4ZmvDoCX1J/XZIEimbKpukjKVt9XMlWu98GN
BA+7Qam2HTkpLFGSecDNScYnDOom+vVd4DvJ6vg5/efKhL6ZKVv7Lr0dWVI4AMAHKsd9XCmFwwZo
PC7u3JqolbOVfBPpihwCyI+1ViohhYnBKGSpuWIE/iegl/r9Mkcb7IlResCyyNS3sLXGkAZTx3J4
5HEkQ6TB+aPaY9gs+Majs3d4PrvSOnUH/RffTYfCaJov8TlsiymClZkxg38t/1TgO2CH1xhrdNex
ZdWDQDWE4DdNYALndzHSlfIJAyf0Qz3QDLQFBipg7vXaCNgZMSPTVYRJkuZGE7ASqmLsmAYNy8bP
fX19klTxf3/DOFDVE6NlXg2k0Wl7WqDE6Iiavw/fCSUHrkNEtoL46UcD3CG8ZXNjljpZJnPWqmEM
8OXkVUJG0o46gw6MTn4VTEkQrQ+267ALJ7MfIxckZQ/35trZAVCZQDgAJlwXAjFyoxRjheIwsi2z
v4LqMcw6ywMiVYBEkeIugpz1X1GQsLrk/1jOJRFEe4oMYK0ZR+a1BNmhLfdlWVLZXc+TswLqMuim
KSu23Swyao886x3c+vIgvGIZXj+m+buQsxeEUYnzMvpZnC8tphEdYwNlO+ilzJu5edhcI3NrCqRi
AeiRLtUlcvBXsGPFntZ1m6/C6CutvqmWNwHVN+e3j2VkT05eCVGKmaI0CqPQqiAp/UskMKH4WsJf
/xVkUop4NlGqavAuAJBY76PY3RelT6OVTb5Z8YXCVDfyQ2jzypN47+tFivZt02pSxcRiS5/QXluW
YH0uanrNCX4tUSbvdbf9OuhAxwc9XujnjbLS44lSRq9COqVrdenqh9allpKVPdO7iiAhEFIp6vJ4
TKwp9XLHB8E2itUOXg9YvZtXkqj+9hw6QxmK8r+rG54S7zuv8zk3lVPPaWILE9GYOcN9TAXe84bh
edWEfSfGfHNMoSolWyf+fsJzxaoovvSOu+cp6OHMrd9JIMiBmBFWTCZt3yxc5NuC3Rjyvpx0clBV
Jrhk+P0xgapD2usQJOEM2gNsIz9Yv3QE4ZSft1nYJqOIKrkfaJuAHKNTYgBZxjQnDIe4gP2PgGfo
ZOSLFX2Zb0tBiQ6QFqjQDb2P5PIB+DpQA4YvsGd7gkAXfbGFxrByfUq43teg1O4KPDB6KiYgtMmh
y2VWKLIiTqXeVG/MwHndLfJiC01haWMYLr0xl1nvpM63LFp276K+cx/+fdVfue0u4bGrXPBv9Ex5
QbYhO0SbtEBxU7FF6crza33jRYAtB1H0+crXGW9D4kgHPPNp3jAtUlEgjC/rcIeIS+kw2d9Mv6nI
IWt6cP1LWVK9RXywoElovXTLH7iVQSWjRF2xd8gDfuQ0Ag7S0JyQij9X05ATDVDOYAVNeQvubyJk
RZWRBsiASmEeQ5fTIunZ+xLIkB3CJwg0JhCPPeaOUhzydx5PHpmu8hN7ZbVtf0ZKSbK7XFzNToAD
V/0bH6tMWiAVQS9tjk1PGCo09O8aDf6xbVr+xNkitgw0c5FkkSSozzEeKhPqgTAM88WLR/pT4RtO
wsCSq1WI5EJdQVXYjz/JNUV3Mhaq0Bg0J1+Mr5jyJ5HzxsXEX+FD0oe+gCi2Cggk9GjAfYrGEH2Z
6JYWob8/1Sche6ioJUrgBUZJck4adopqobEerW4hG4/Ul5bks1IwXT9lyPk4/t0+JR7CgrDVFQ96
s8tLPY4tLseXZN3u8j9ccG6+zheaJat+IL2tNv1BHuoi+VI+SY/fZSPxDsQej0GkXEM2qAI77Feh
B0vIXe/dKog9E8OwPu28Kxvlo9LcZi3jkk0vTPIxOaGoDYyJgMfCkbLjOKzZ5HYAUxmCOdQz1nzU
ChtPt6srNXQZztuqDGBbWgCiv8UiJ1rcZfIC6UpTVVUE8yjdWiaQ8wF4O5nH0RPwRq3KYjiBfPi9
qTOr/Gz2vXN3bPV2TvCvqe/hxnoPH6j7ku3amOJX5YOynjxFhzPEH9cmpoIebsuU9WRYO62FsD4t
6+z52BNAG+P9XjkPjkPxIDXBQF315gtnpHRPHuEdq1U8Kqf9g5bu13JY7lFCG2YxZDK0p5q3n6QF
F//xLJgAzcgpfIAQyr6h78bJkomIEbIAjfI+SkxLYKtoDFytofowvXMoP4/WpCHX0zpXyKg3XToJ
d+ogqNQY1tf27rDk/gooTsi81Ev5xbJNYtTChiEr4KGbwOTInWIxf2pjry26O6Gxmx/3+OBk+YLx
hnqhEJrOx0ofnLcrculP+37q8S7ctoaE934SWFpqDTIbJfXFzFm3k3q4gIU46bSqK4h8uHLv43pB
RK/cDJ7PRbL75ZrBnRfY91zAHLDYpqLfSOTHWTIBpLWmR3Boe22x1ihO1OC+dH6vLf+JJtC//bN4
P2GUz/kPdg+lPKFxRtSNyDlEyUs+5PA6OIHXj0E8gvCfiiMD6FWXHyNluz8ralykgxHj+M5HLwlW
QH+cBmRY90QN962zLd/+k42LPGM1hXa0FlcqWT0z1m+8uy49PL9NDsyzIaPUg3iLb+gPzegyTkht
jZRqBsdrLc2oNR+4Cp60AeZhOA+Kl2YMDEE/QmHAskQ63cPItsZ2umMA3Ph7DGA/TNl/sRUv7DHo
Y2d++6tVxMu1NaFpj+2xJsL3AdQhvEzrKxMIaRDY9wAJ+7Idsv6fYqXKgzkIz3+bHsXJH5BkyNrG
EK0CC7jnzFLNGOJGhphZDhZ1P7aSsG/pbE/qDZr5zHUNoRBFfbYCFWYezqBXMrixTHRDXN+ZyDcV
jxEwP+BrlbhFuLvS35NmR4clS2/boIfJtneANlwinUQe6cTSwgS8ga6zFhR01VzbBwnOXUK3uSIN
T0NYOfr9BQPSWRzr2sOQAHaGRR+pezAfsBAp2QkVLEyi1h23ibRU23X8IhK2LNucmiyS6EV2GfQS
IKOVLWoHD3Dv1igGfpt7V4dTJ3vKTxHjfR/snIuGT9x0i54W8pXItElV4ZUu0nh+9Wxm6Ws7Zad8
jVnIYazA0f9tdm0wloE3i4IHyWWKjRm0iNnaZD7JFT1K7SJFytNUMs5zEx2/cY+BA0ARw4t8wIx6
cF4x808YGmbKT0hrTUopqn4DGXVH3S/tGX3SknigWmLXj4AHJsXczuPiF1FrUrCnVLGdULBU1Ez2
UdpMQsAR3PrFHbrgt4mNdRNrLwrlKhAfEHzMWo/QrtxBaKWWu+wSnCrMGCXhJnanlLbBGHaFpXnT
yRIvXbWhCUu2YYPMJlilF/Jrk0I6MYzjZVoRoQXJ3BNlhhbv+LPQCTSq3tfJQSWRsTE/WQPQkWy0
IQbE/ANDAgCouTCgF3LWvzip9MPHVWhIbUae2Yc4585Nd2q3QLJ+pEsyxQ/1YYLCNc12xccaPMYy
iA1s/S9B8BQX+E7vZUdchiBb3RkP6WoQXZWeLneJGsWoCw0eQhFRMBC+vXqr74EOJrA0aXF/HeOV
DRYF3fYgSsnPI1d3D2pbIUksAXkNgDLpqrhuez/x+6BEjcygHMWtuYUuzVICgyuUTSLI4Zfwk4++
XiBlNR0ErnXLOGY8NrrkbzuPnDAoqXhr4vkcJvcu406+mGjjRwvpIcA3ar8DXSoIWWB7cJEIjS2k
5GJEXJEEr7DkcytHauyiQNj9acFCE/oktBRTXoOVjMqAeI3+Z4Vs4U69FEir4kMaWkNToqdfr8px
uR9XWnCGpJvMTdEukaS56/xOvNeY2D0a6v/b90cyok0BhIr0KImTSDR6uujwkD9UrfUxT4RZ5xDu
YeRLqew7BXGUmUSCy84HwCSpoAlFnSbRrtWf0EBJBlQywM2E7cMquhZav0JWArpxYx1mSAw0M0sK
I0zjZVErHlYRG35fr2sGykS3COnS2ZMeyjgWtcjqCACpvUfmFlsIL5LBWEWwGV3wEmaSwpB0pJ1Q
heSqNFigUCBC8Ati/tRdvF1y564dRkBMHIEs0ygkX+KBzVEM5uyjlD53cjyAnwKZDrEMdBfiRsi7
/YHXI2nO3h+sbquY33Y8iyayLkwE6vaTkcyVy6cH80iO562WKjCXV4x3UX/A18onPJ9dH9MtNbbh
p7MW1MtU6rzvNcxtk+QEOF/cJTI3MMKhV+BCABJITJpVQ3CxpBc+/4ebNWD+/2No1lAFY2eMOHzE
248pR+ZPF/dKWXFMVB9dLcqA4MJupwn/Qiqj9A+SNGk42pNPUfRCdWsvYJ/xLzRT2UxG1K1puavS
cFkq2BxieXr0goAt60R37jY1JCpLs8ZeHSMG4skpW+/1PQdGilgPKYQr7FzCGsUF3VJCiLtCBjH4
9s9ZL2HfOICxvm3r1bc8zcUnHdkldKiEPpdk0bHg+AReMlnPayeWJvR/GXjSkMxd40o0DQNIRgdD
vl4BevwXgxvJTghbX3o5e+f6eY2Y39ggT5UQ5scZd2zWHz9FB3pljj26KwOIC+hDzh9ITkBMacs/
uQpYDiTRymYNN8qZ4OAxwG8suHPNR6u1Dqp6oRFtHN+016bQFZql3c6np8SjnCqaJqco6LHVwA1N
AXPzZQmW+R1UodKWBVzr4wxYOWuKqfj7cSpoZuTw8/MU1+41fN6uViUaxCY1kuBTpQGKdq4MY+KU
wDjj7ycx4CbwPiusOnHgg3WDEkzqfwonE45ypZ5bxnhCVw8p3yjGcgKhyvQi+5D80p2Fnz8AIkqm
+FcjHkqLNoenMlygDQJLaqHoGF/bPPSu8cU1hiezAbTNgJ4WxZb1mJ+5CB+13ae89hJz8HrXI0SP
TE2L4eN7AjOkXbsmLscv64XRY31Co2/O/B24kYYv7CZ4bvKwkInfQ8ChkmVV0qcJCbh4F93QtgY0
1omFNMjjHi8yPV+vLLvyffnjPAOub+eNB63vwWzz592FBo5YTIOAl9l90mFgFhJl1NUpfU3DRk5g
Y8/78DmG7c+8lwt7tEBeGQI5HWPvZFshIj9+q3A0l2wS2V6k+DSwbzt3E39bZK/cJDoinFm/vUDU
V+5BHyOGfX+vciboWD+4K/eAzPkRlWZu7fQkSfNCIVVB5S4U9b04bVJpGm7Wwg0HtZVkGA+7e+Nw
W28QsvmrtZJpCigGOGzoIU4jfC+4QvkCLTlgy1gbl4pZeFMCC1wklTrQpkjhkXOuinEPB3tcCrJH
V61yw+3zga9b4I+BXMOoNYjkwA8MPeA3CQiZl0FRld24yYuG6nw8wG98W2ULHhVfg/A0HTxDtbQQ
n8RNL9wCUE6C1JhhlUkYz+klM3Y1/avSCF3JQr/PQBnRgkAkJ+guUlag4PYNcp3Dq0pCE9wpWezt
yK7vUljA1TqHgeQkwXvGEGFNtyLaPPqk9DgQC3fmsV28+i0rjhK39BEyyGiEQPe5WVn7m1dVTj+E
tKOT54eOesZQNVcGKHpurVycxZ+G4BA97UpeJ5vuNgqB9BXvUpoc7YRiR1B/Wv3/VPJNUCDiARUP
ZdMcVm6AMSwV0KvoEYHSvZC5PySbRNvZhsGZ9WfPOXDURgQEQGXFbSCszSCiq6hWZ6pyGn8wpoD7
Z/EI4EyHZ1KSwIyk7rA9tYQkggrsFl7k9DSVDtjX3vbUnjNUG2qZhEarT4NCQdjmZoo8eMwMYqet
0J+224xl+by+A9p9VaAL1amq9xuhI2FILO7qiQIgbztE1R8VnU8JYRaOrSUix2yM8YTPn4AbFs44
XRvKPCJ6OcrOOoEd6+YzbPREZal0vpKFMha+oX5gnLtfk1I40Q+oztlJO3g/Q/hNvJXE64M0sONx
ZD1u58/G+9DDLV7BMveEBEAd19u4Tti82kG0Y4EjQRdYg7yrdl3hCjbMFIreSPcJfC4dVeU/WVhL
rA7sZtAWTh8lFT0LsKosB7iTiBAYdPvlEMM4m+deKLkJbrGsGTPbuMYn3ILEgJBAWy1IWMK90Gqz
PI6S4huYoiKGXFYOtzFA2VnxcQEMcrGuVjdnneO5//NYXurk6KeMm/I9Js/Qt7dv41PevTBENtmb
wlQZmGzaJ0m/3XA3MB4rHbnmXdCgE9RJHRRNWOzZsV/RnjiNtZdwcCdIHLUVg0WZkUGP4/jZGTi+
2KiJKcxAt487zM3yQ8WbDKxP11PXKdYcf1tQLc3qYyPQG7LbWZE6+ZvYtjGzPtO+5Zmic87U3lQj
/0fN+4DbE6NXBoZiMl2MsU7br+yxlC7r5qkJ5Qdt0LfhoUEp+S0XY0/JKQhx77FKK2r/PWX6C3uH
DTand+mazhDcQD0hWJvrp9hiKuk5PTpw2jhYOj3AlmAI/GUGRiB7gklMOmkLbwM+VUoqNxFGrUBb
7Dnb5xRfxI/XPJz5t/quU173de6d8cbQVeGL5Pl31eP0l6/CmdI4m3rkPccORzv/Q30Y+XtJj+0B
T1A9kQlxrEppHCifU7r5XaSaVUXmadveFXPmMP8kgzLh6IuZTVklM+eS1amHiO/lp2eTRE7ekfpR
/ho0jkXMf6GhLEecJMhXgUj1ZqkUnIBEJpNIKtahHHj4oTRR36DVUyAoqik4Meqmc68K0goOF+ot
gUpyvkFicTugwL6hOmWl2/3nxe+3EWwzlnvTiFpxLkp/I0JUVwqoUsP9O3cb9dE8VUZFF1mO3adU
IIEogEvS2lwLSepDOLOuuInQWtOqX5Vaa+bT+jbVYiVJvrr9xQugbujNCeP+2oyFflKiCe0F2eet
z7Jl9iraPCqr2+dXib8rG0kk7F2JcOZnGKwBc6IunhIYBGULQOJIykv95qAZZzI5Lks+brshqGQb
2N2NzLHN2JUgabkH3arWvCEPxNLYr1DFMvgqFQ9c1r7cJdhHPG1Sv/6Li2oXLUGU2Vxfgd5+PCgU
RrJJ341zXj6aLn9rlNluLOtaXBxNI/OaEY8HB71bsbj6AY+g6R0NNUBLvTFgpQ3uEcjFFueYF5C5
PU2xRrJ8GqzIbw+1yqozWrl24bEpFOpPu6hXhlgr2jrbPtG7cFvR5ZemBmbQ3MgS0B02qN8pywx6
sTIqfytMJw9LmN96Pho7gDqiAACFU8NwcBVihmOCzTF3H3ys2IuOa84Yy5oUSW/+yqWLVTJiMyXl
kefg+3xaxvvZSNZ3uZggsHnOy9V1nPsbOGkqpC8ZWsWv259Kjn516LdJZOmT5eABsdpc/A80ECMh
u30s4TGOZQv+RyJEdRWACW3n7mhZfL9pTNbFSvPafrTlHDaMbqrTve+pVz8KE5AjChdQoJs9ee5P
ADo0HkWCTF3hpCOoIZRPwarLDU0PTpCAkdkBiPFCde6NyS7TLjAQohyS/jWvv4hLS28EIOXombPd
lovuayY7ReTZsFlP4Czp/SZP5ZBPJ8HZgTN7T84PqKcmIgpgumbkDRwYyErD7WXeT8o8sN9QJue3
h5v3a7KRxcnhWNJMmfR+1vR1LoGbTYT5zKbZ2rh3eD549Y1I10AIRihJyXzbLpd90GcrO+m1Ekmp
YJ0vboWGj3fpxJtrzWs3zBqO3n6ccUw9fbcBerL0Ru7417jcD+16z4uaN9DiSkrjj3xaoYXYypXt
rAr0ijXBf3eyRpbMi263vQ+KG5vwHuTq2o7DrjmnRFlpMySJhMwIpcgPG7zZh7iTUPdAAsL2akIJ
UVZrzZEbgOYDKY7PkJW/icE3JwlZqd+n4MpOz+Gro3KFbRNBokbMyYbT7wejB/zKyoTd1BNle6T0
o3keb/rZ13fLgcEIFoo0U75MlUFFHyC9arFW0TFEINQGfz2yBvZepP/7s2NgchU1tAe0cSAtXQu3
4iEYTH9OsoBDbUfP4IX40nk1zj62gJCEnJb5beM4On+Gs30o0Pg/N9t93FbAdQ4+N0MpxFuHVkMT
LnDsWZ7lhGNJ6o76f6kjUVp5ih1a72aXVUYkSM6iCwHPjSznjI8r8tbn5oLqxvBOwlxstueo4m0x
RctHNL7reLoKb4Be/YJCzoE8GqlspspivPSFyyIdFVy3ehdmZwLtbcSl+h6CXhDjnMGKD9mSeInx
ZNrD5A8NWEpZi5VNxXd3YdlXtxx4ki22tGQvtlM59fO2zSqZdjAFw2y6kSS0Xz1cIWFYleSOuBur
IWY8VbL+bhOeOcgRxNYDe7igj+TrN+g+lVFhIHwsNB0RO7vhkiPfvZ1Yt2t+xtt5c2DtcBbh6oNA
9tjJ63/ezkIVIexvBv14nk+sq8PvGFYBXQ0xgxI8pHTg9TihnDxrW6slQbLJrUJXXligJPAs3jd8
ksDiGzBceniqe2CmBY+YiF4bl8sCsgGBfTkpEQCGLuHnN65m3ER2pngBn2kK50hS6hSeuqbAKxLg
bfmjZEHwFYGpI0MfRcLJqd+Uu7FQUji/fic1klXG1HwpJSwWHeYj52VlqQexX7hiqAMhQ0qy+bGa
TbGG96SGipfl8zgkjvMUXr5UhvLEZpstMHzNFF0qMUGjsPFAVy1WDLFYz+BNVmyt4rsfPeBqKNdF
cV7Cw8/rT2VA2KMLeLyGDOJYgzY6xc36qj3N0tHk2G6ZVG6aRfVwKewu2dGFW51ykLVAKxGj9gRG
+Io36uAxlsgMkGjaaaalkce63ZpSiEyvEiAwzQf3fCwYEe6tP0GN/SypjHAiBl+jQ2Iv11K8FHls
93ddTqUqfp+6QGlsmyT5hba1ivyrMuaUKGe/ias3JFQhThxF10xgojlLaKawT5OPg3hj3C7n4UIp
kWj2QAJ9kRlwHutCX80uHMe8VLABxm5b0mUxBYVrSERh3C+pzZbHE1V2VIDMhblkOPTPgeGOut7S
ZEw+G3wrNB/mbxaXELv8IMQm6fFvMWqZZHJRMeb2T4frMNV5AcPDjOAicYaIZQrh6AJ4fCfFhDkx
Je6TXR8dJ4zAaepMdlWKJNRW3+OA0P2TQxGwvKXxCV/YsU60yKry/KLLcK/X3M7dGb+tm2V+Yi+7
0OGoAP2Oew8hvID51v4fTXDB9AS3hpENf70jLPjDHzyWKzjXMIORVguVqjiyPqwZJLAbnsfxY8ee
LLOvFXLgLg5N3V8R2rp6AxplCnPp8joqYFIDHWOPrq5LN4HHoMTymyr02AppwnZ04z4YBz3bq6dz
UwU9vcBd9Z+CvJum45vl3Z7/e9r3M6XjCuwdyikzTLRho93pztrI4jS8sFH0/eyKbgvs1uaSiSe3
B5n4ZjiydO5dheX+Mp+5ylJnBus1OE/P70ViNvfDqNSXywk37GF7xqeabUUl31n9ZXztmHQ4rq42
ltfzKkWgLXayYtt/rdH/3O5hxCYzipPQmWkVEtkVHu36V9RkW+XkWebORot0fHCGqshnliQzq0pc
vkQ1mQ7KwSuvtvVNV/Uh5yGxhYsi//ebMCVeHHhEiMzlN+v2BIzUSAnRvhTP3f6RUpczQsEEcYRT
o40pEQ/e+hggiJ+NFmpAgqAW/ICRPCvbeG2j1xSd5mU1JMghVSNohOZjtIcXf0cPrwvR02PWtR4D
SvGtFsIQkA9AqAzixfZxafEpsMJ+EiYLbDUH/JtL2WjRRrU7ItuQGbwPT26IRPrMLGPnok4026Pl
yRMzx0a/IK64Ve9qUuojqmV8S6AjSr7cPJAL5XQnxx9uUwDVAtOSFZfJRRP7wjfVsryC2qhLCjK4
Ol5aIWutYXqIJsZCbD5N16+nbpdMz1sLeADCgt1XyetU85C190PbV597c3ZEZnyukkgfOVblxW3q
PpKLWLVg6kh1sQ+2DbGRIdluDLdWxTk+LNLeMOAddY+8L02JU2RjDu6n9P26NuWdNE/VtVGqzS1+
fXvbKELNrzZLBawBjR17VG4HMDc0YkpemVrywM9xYPHFctEjBmZlZPrIiCr2h1Gudy6qVs0cCV7K
75Ji17TBKdBneD/oZi2f8srZaKDNJN7ktpsUZtjwhwRMR42BQ2Ahk/sprH6XKLLjEKJHtSzrG3V3
HK+ziS4IAa5u2xBCH4MZo43JW8eMM57Eedrna1PDgOPTEwNIWxv0wsQtRtQDidwt8JHnT0VKyAR7
404nzOSHM4g/EklrpembJVfTYrCts6J15C5asknXcUwZFkFT/q87eKQfWYKXEIMpuwbHsgrZo4fs
4/CNB4hlmcPS3Bg5zaG+vaRpcywUm5yN+mH8prkJwFWi1kq4Jq6EeqkktpVOWrXcizSK8inECXgi
QM4+IRwm4YVbZNyKT2ToJiNvXC2+TOl+dTsexssdVJpgHIO561bBSitgJHExP+B9dCoH/XNpoljK
XGSXS7RqVhsVYegG4WEovklXmdjCMIl54i8sn4boWDwNlekLuA+aZR1WZvcPz7YD/p5+O61YojfG
XHVRLaZapZSo2TztrpGgu60n1tQ4QbOpBaaCubO6RZXWzIDxPnypyd0R7aPVL5T0GA6XefHzSksl
+HYI40NS7VKpLWUThtL+f7B+KVueemvN8HIDRqojjpmiLLOGCbAzzdFwIykjLCsc05kclcvifzpt
GZeonc5xikaAIBY1IALOwOln8UNKr0t1ZShDWTnV5FHlDfJTvHFBZxDwVD46z/Zl74Q4FlaWbvzy
eAJAes/YsYlAp2ypRIUHS6tv6I3OasgYl6/hcpZUHvZEcmO7sFnFuIUJjsRjnq6I4VJK6GFyNC6d
xxY+EQHE05W6mmiEWW9akJ7LHSjLZ/OTEzhzoY1o02Iks+MjKVTG10YU8RR7mDGy/ePvIBJ1E/+K
iwAqHxDgG59Jeyszmsxk+8nmWaIXwY3xsGlkBjWsGW7xWRXPXMVtrPFG914n8JRSrko7bcnU8oYo
B9gUPGTbZtb6mtLVta2zwXPoQf6qijmKT6wrgaFuCcz1GhcFI26sOyrL/HmkjhWKyPDjj+MPsE3O
Yzd4htqBGvjW1TheMGKQfkS9pwKWGSLdwlLPY76fAxZZjRASflmwj5Le48aner7LwpsQyjCF+NRF
GIfXiDZgC1/yZMwCq+lF5XIdQ5GgG3t6pL6EWKMBErIV5fVkplVpg948wJup/osZUXRVUCVTqyIr
LMK0d9Is4jfnDJdmgkRlDJgwA9LAONQ2gniDuo6AT8WoRIBUM/KE69K6UsbzJuA0ll/DG57RRxwz
1Scxgj7Ih9ZrA/jIr3CGo0mnsyuuN1v2568pc/mdx3EMeCVPGUUS3vu8xjP1fi3mB7xO6CVVD59Y
2jxJ54ZqMaedQGDYjZMSUVbiwkZXBjA8t7R1HLlRcq95xdCl4+PO2hcMS9hB0ox13rnGzFL5HmaF
o4bt/Y/FsPRnvI5vC80ohVBJW7lhn19uc43dokCU6A7Qh3m69dZZv9RcX8cFJiTi35BSanmt3oOd
W6QwATwTN817AK+TnrqoE1Uvyo65BQF+t2jAF4xLKUO30yyL6wgjL7S6l8AqAXg6abXcopNzk3z2
ExFT5qsCH5YSiHRLQXAObqxK0WQx0v4E9lLNGSfST3WiSh4IG94IwyYfIFLdWmrlIGBuO8XAq0Sa
DK2t9e/hR0X7I7URu8edTCXtmguHmtG3CjckjJ5JR0nRAZyzK8pmUOr/LthoVZAGkOaiIDJ1yNMF
/wQST/ocsU+uguJktObWPqhd09ReXIK12cqNE1ew5V81QRsj+5jk7L2K/Kd2H6vO5/SwwWDuacd6
MzloblwDdxZCKhXX/FS6L8ofFFlnvyCzqWIYssKMOLtoAtJ19W6omU/ILByPG0GfJeil910eRAxn
ir82XgVXYbi9B0TD78QrcXWTj1KIw9y3ub78ZUFSNj7/VZ3/Q0LAAhFRA3/xxmoB35O2gCsbJLLd
TPZgQOj5E4Dg8zeAHiANi6dr3ZJ8a8TPEGCxUfD0Qd425eOlaIGLPghBzDpFxocFjZ48mUIWJ4Xr
wYuNIbAyfn0nussGzvtQhRO0lDxznW73SpHRqYD4K24TIJ0QLR6dKCDB8GYdFt7slvAwTplISrWE
FXZY+XLV10HWwLfriJrKYyeqb5RCub7XyATwS+we1h20BLowP7nEKxXyJrQjYf2rFPZmadoC3jJb
zFU1kStNGisScehXLqpgay7+KP+yDlDIfeR5Bi+96Y9JRpNx12cbvAvnmZHEy/2eQVQ5uvqoDkts
s5MplVO3JrGzkPgpT75qiI7Fgezzdya4idLYvM9MEa3zSk/Sw/4n1izd2TQ1NgrUZH0004g/JdHm
8FlYFgTGBZ32m6Cmj5pP2jSM5GFRXV4s7ajZYPzRbPxu3JL9tsdEQeEMKzBQ1Lrp2fHH+tB9i+xb
g/Cfobc24dKbvuxbDJjTL8dLQBIC3oc6jj5M/FAd4Bi2K6xd/uQQsmUSYIbiZIm1eYOO0fmHVvrI
8ZYu1YJNkSGH4Fwti2LQ4Pl5/wKI05Sr/rh2ZoZVPGknrLlMCVE5hN42rUyTdTEMceyiZmwls1Zm
e7DdWycjjF7KaGUSKK9Z5QJqSV7JSaVK9rOpjZNx7N8PRwK3x6X/bvP0cBjDyp046NbFcTchzlZT
G7E4sxFfo/+EPAthpho9JU+NQYtmV+mqU9yBKbNMEtgSeZsJs/fbKA66lMAhibO3eZ+SLQrh82gt
jP6D08C6VBJDk6FYk7wr9uN+2NgRKHYwlfWoS+b0RXLpz38gfIgTfb3In6WyqFAtFRZtC+I7B1h/
JueawDMwDl7/DotPrFuAg/0+JaR5t5SOInyGIkhecw1cAggNkzNgE6KUY1AWPax+UY31cu+Bqz1s
C02h1gJD0Du4TNvo3foGhKD3gtoEl0OOToZBOyS+0Hq0ZF8RLLrX20+oVijYd8lw0n5XSfgSYdR2
vKKQpYEyH4VFbWH2U1fsspMYIl5+B7gFL5vdxsGF3G+/bpzaITAgfQ4mJrh0rM6xrw6RGNBsJM+y
VQJ7C0ortaXrF6Nrf7Mi0ZmluWssKs8uvWYVJ281C0M7TVAaUxobR/hrLeqRJu5drVP6iPol8bh4
NEQs8liYyfg9rKCFZHkRckLqM+UOSnT102SbcBod/n+pAA97uO/PHfRbtZmw7He3lozapcIRVC0Z
MYGXoeqUgOcGNNYMLNWDSSO1+/fXfjnekCnSc6/D4WnANHBbrLjA1rPqHJE9VNY/Gp+0bpgVA7HB
uHQcjvuaz2TRDvzhEVciBf1Iv47UZIwh/eAsDSLHp9h5JLr0lwxwLl2+ee7bZsedGN3D/91hjtoO
0IqGZbCmOGzE19XVlJO137ukxIL/l/tGXcZY3Fqaj2ikzAn0z5xkTEZ5GUAw/5w5LF7UHD09pS4r
zcOTnhMh75iensRUnMi3eUEJKgLtnypy1TkND6RWW5woYyqjkyDi1gMg1RwE5SnwA3fb8CRXSDVs
z+X7tEgvZVKsd27jgkO7CA3zUgjUMNcgRiRdQtrtfC9a9ioTn7hMjFLmCxWxRfyLcyHFYCKVy3MX
jg7ssZr1vMHNQhMJ13kLnZinKP2Ql4aSA/fYPu1QLsAK1kR9A+KqA86KVxPANm8amrpoRo+AACh5
nCItBrJdORwP+DDE6f9KRyIAuIZMiYSqZ4wZsBsL2sJbA7GLDmQbJMgiis09GE4+s7qd40l/RTUF
57yMbjlSNYXJ8tvuNwEyX1jYEmSn0dF977ALQImldBvxDzNHHNId29z90mAh84PW+1y5FkvAoiG3
R6S8dPBC5gkScjEJIhZSbvCYvwXkKhdtPF4YpXNyvh8QPAtGFulJZkKNuqiAIut0v3Sj9zC8vCaW
7nacnF+5ebpt6/bL0LTlrJILpdAcwKaqJFY1r3V1TbD5QePvR8ZMk8f86OYThbgMVk/Ea3Roc7qQ
6uop5urK8IphzCKINACWwWCiEtHX+xeT/o+JAcM6jEzFGu7p2MxvLGjyLy0I5nJaT2SeMm3eA2bo
sY35VXO0vehohUuvDqIW/O1CnLUgyakfFGU5QnG5nv/SahQEhOuqX8mwfkyreVOsJs4senFril+G
EWNMPT2FtI71obx0c1jlw6NWLO66TiCky8IC/NyQ44wWN5X11ZnAxLxxjwIyrWYN3ZhDt+vWIjg2
CGdqERP61uP6RA+ubXXxC7fPH6Qd0cliA4j9/jJviVHKaLvT0prSQBCB1qoE6Rl/1mdjd6XJ9pbu
3PPf+uPINZreTSjqYpKTcUojXjL8B9Ip0kKBnVf7KIplIVKuX/V1ebCKB5OWNwrpIVIrFQ0drt9i
RS+9lCTG+OCAfLW4DyBOtziEWp/3NpAwRPTZxwjziBq7v/kolodyyejtmj8N9fuk+1HsTuRkcr1V
BQPQw05+JCMxQlmdYp9sAB7KWMhW7babl05E5GhuaeFIGGdUu0GVilMKJEQV5ygfNS69lnK3kQwQ
/xakLpZsPpHwWNPylE+xmPwGdCxBe2x16Iu5o14isKk0iSHwJWrA8zY3HbnFFacrZT7k27gYTkL8
8EwYkrNMrY5w5hDLhB5cEt4ColsV+jRcA/cXKRIXW11GHnQSg0LNa5vdifBI3FUNSkt/JYniTLTp
Tscq3TjouLHqzREVC2gTi4gP9G59h4CDWeonmgsPi80/tyQQBi5kE9FxlVHXrZEqzDgP2cho54IX
zyoG3jGV9g9vCXeSlTE3RntcqyQQLM5V8FdpgmJ8HItrQK18tYBPaVjrFIbk62PTvr8JpSaxIraW
Dqt6BN8P4xK+dmguGqi1t/kI67+GaHM2jdSyz6UTVH3IJQWN3O8w3CBHyj/boY8fFqbn9Njvl7R4
2BC0zMOzZ3YyZEef8IboJAudtp3aHC303hEnin+f8jZ6F6/OzxXGcCdaeD0KPzoSiQPEgoUzZfvn
9aG9m7EWtbO9WtyvP5GhSNrcBVus0u3D0pvzCqtQeBo29EV5abivndSTvbyynKywY0pLsKqcBl2w
ejBCbzCX3FAp6FnTVT4l1zD7aUWyytEmU7c/pLdSXZx6LxUjyzoaoisN1upho3zWf6OMRo6Jz9Mw
4ZLbS9pjd/kurns2FQJV6hxvt/qJGasm3qEZWrg5J1EgDGJG9wacW2uCTQiDuo32M43Lt+0pL7kJ
tSV3NOWfxDYCakf3QpWC6nlzsLnx+pRyTBEaplq8v9NlAZnxO1wHuGwbrlyXgkQjmws8LKzeAJtf
dPfPI9euaBp1TfXPg/dYkpPl055iVRcnoLGg/ljeecTnXCSW6CJ/JEvn5qROg41CM5UOiou1vNAu
ttaO6wv2kNtOvzTPWosSsuD1jxRqV7AEtb7bZQbtEG41kriF86o7aDaUt2fpYXCY9KhlXKZZWj39
Rg4m55HbRQyELHhVAULVQJj7QjL78uh0DnM8bkyMHGV+EBxQf6pzxRXnh/5kgbgF1WocSLHhNSq6
6oapJ1wDr6TipYuOZJ9uljLN2hZNkXrZpS0LrWOHXVn7tHm/hoFnzSsEoRQggdEyp31tpFwwmyEc
fZgJLDaSJmNB7KThFCDhpcuHJXNtmitf0cQ3SAvkQepyKoUdVxbdhfZvt9LXdRfjQCFDfH/MWpz7
yIdZwfAsYO9J8OmnDECcY5TY+vgphvhEQclYPPTDv/7fihZu9QVzMeGcHUyMxZuvqTBcFWpesn5M
IMYByswnGIlMXpQv2HySZbZFcd4s8S0lZEUEkP2V+iLtwt1w8MRFZKmKLphF6K2d2dGA6PT+dWNf
Qb28VvH4OXcNYdfNVs7SJjU6Ud1uFB81K3mZIdbIGJ9dIiEW7CLXi3Uz3lbY1qLZqdgmtdu4HAXG
J5T+6PDzvlQrFwn3rQgifjdaI2jPjn0u98SHvaztcu1Nv8sO/g1ykwUAMHIXrZEvQ3kNZP36XdoT
FI1LYvIhtJKaozGZEiTiWGUzV8p5pCrM1azK0MV0Y/OZBCMR/vBqJirbh61WrsMRZSnecxhVaYlX
f0WzpTZtxEFyegv0jOWLoYpQSgC+mh8CjY9qsBT/BDQcDM+0+PyHF1zEJtioWtvE+XzJ/pWJGxS4
gebL/j06V0wIl29mL2zW2CSU72K2L3NrweF+fymv5k1EUUEdnTTemE05K4Ei+NAepY0N4XkTlnqC
vE2PsKWiG5nY2SGDinLXTHQRPzb7GN7UXc3p8Vwb6b7ZsKjfCMavDx7SS+2bZqA2cYXcCBdWQUQl
QfTcUbYusdK8xsb9d4UqLLIou0ltQGHGZybCwdXPqB+Twh7I2fZ0/Qdn9NBVOUxU1rwLfG3jjZA2
WQH2sIOROYs6isEy928zGcV/xL1h1sRyIXLJJ1cNjAjOgvqXfDbUfTLrWvtRNd+zkghQzXjTTRz3
bwj6g0Fph7FmnxjOkBN6rXpUeXU3xLUCaIal9/5nRmO4Mx6aoiEObSNBiUokRmYIJi2XlrDz5ruz
Db3ajry0th8of7E5y8lNQZMwldtJ8+RsOGt3PSHfeebkC2NGzAql7Eg4x6C4ik0SgWm6xAfXgfjg
8sHLH+wnyhp1+d0g605iufIh6mfr502fH5RWbKmH8OhTlhjaBclDk47+wCXMcpQIPsWKCErClDM/
Hx55cVgzvVyaPpVJ4gpo7sG+jbOMQNVNq/v5FQxO0Pvak9a8n/LMSGVrTJkLnjBeZO3+TXns98GB
Fo2ZRHWdEbtBTijF+bN7+XvcgP0KRyGOH+o7QXxWDttV5fD5NuQYGx9qJaLD8pnBlscvyIy6PzxX
nEwdWL8G1DHqi78i4ErbLu+eHeCi2c9MhZJ2vId3mCJYxuDgnnLcJvil2e0Twi6M1QP5GASw8PMV
Jl+B5h+ZZhaqWTFha4WrTZ6nMYM7d6qF62Wg/mz/UI+EH7GXxdDMnMMOHwhfTFvG5msMXCHqXPfD
uVb6LWg5XQNV6kygGP/jckaPagjT06K1TnVXCbkqwDE+8S95h49D9JyRSXC7d0MChQr4rVaG2N8t
v/iX3lj3ZjFO0SWN0D3xPILndHLKI3q9xIRg02fH9KMfZ1351gBjzChniMJrZwn0jpYzUy2YILrY
EjM3ZeIT2e7fxcgv5D/Ffisa+WzxZ3e+/fXZeLnCocXHst0qUBWpp2/BkBavj98PNOnOkKAHrcAL
KW+1NYNv81YdJspGt931PqLEDfSdMZihEldZue/AkWoj4FKxEjrRoKRrzj18O/RniMNjE9EN/o4B
VHyWCVVnzV13+hOE5B/5uotM/fkXbWX/Qpzs8CIz1o55fyK5paW1t7aehVNNowJJkZpUCUPFQRXb
6IgHNaGWkylX2yXZrWYbAq12HTbPi7rxtNsm7mL6vE/idoPVLSvMHnnU7fS8UYbUhO/vrrh6sOCz
KZO1t1sxJHChjk97QRJA0evysalyCGy72ZwJTJ2TCfgVqgdxDCD4ZoLc96SQvnsuO7xgX5LY0Orf
YOPSE6jxSJjxUUlCqz++BVPsllc/E1IOTnbKYWBRBMhosc5Q5Ps/h4vFpdFNvbl1Afh3bEdp3G95
5kZdnq7MsnVb/4Ujyzco0E1KY9L9LFEFhbabQ34X4TqziDW+Wsy/xt9F/U/mvTaywC+LeHhsGtKP
/8zbf10LXTm6+qH22UxeTTjzp79J3D29b//St91+c7IvpNoG5Vq+QiMmtGBBkATQKDiNhUaNnZxy
H3HwrxnJsIymVxtWq+71lNbw6oKhi7aC2DKyWNlbRJxBpHnw/IHewaPaSpNajcivEB+397bumIB7
eA47XoB1D0eMyXq0BKlcmoDtPmwSZNUErYdv3E6kGdzioueseD3aIz4/Vi98lKy2Ss9enHE5Qxsb
m4lQ3k+tlBsDzovbIdVGQRiveB/kXet0chkwe6KQUm1e0VTVnr1owyFx3CHXx0DlcYjv4NCPPn1e
KofjHCaCrs7RIrKP+nHfu2L7JgwNdtL6sgmpqmdkl4mcVgkiN9TpOWVkn6IPaVWHLgzOI0lSSAf2
h0xtTlXsoL62G6I7IIJXNXW4F4UsJqRuHdpXn5bceUle+wl4UgmQ8YKJ4gjtraCROcVWBK3duViR
nbl8Q/+4MYFyR1943Dz76CCPz+nt0ezy8h2NuLiVaMU4kMAOBCvxvvQh0tdS//SkxVHMraASapt0
Y5BUJbG3RJ6GyBiKhcu3dVhiAM7zEOWQCx7yQfvLlCZRFCXA8a662nBHRoReRmg/0hnPm8kBfpRm
Mu6nPfoOmuTmvmEBQC5gl4Xpx44W3+uT5O4C5vJQfmrAtZIHtg6Ov6hThEbayBoksAZyB/m1I5GL
SCpjFafXBRzgG1GEzReudiOYD6mkRaAED6u6aQBNP2kocDfgRJXjurOIsY6HEElu+QrqYRqrrxU/
vq394zaSKT7b6KtE/1ll5um1Hm0TlDMhzQXnvMc+Z4QvqzoGGVRwXxn9Kn/VV5ROpfjtZM0KR6ix
8bGYV74CkbvEBFlsBUN9l5ulXp7dIFwJaE8+hWVyiZ0F3EKS3HqDlS0dGkXr0vVusE9p+WYKlY1a
BCBgkqmVnOi2JTbC9clWXnsiQ3JxojGFfnhwPByOAjUZEo0k7fbRoYrbvWCZ21PfTJ5lWnh9nTyS
4vJeyV6Qvic45RYZlmxQrG7glrZEeuqTC9OmGLmD1RgtKq8XQTmponMvz/ypkU/aklB7WDAoTwAu
PXs0jc4Op1O6QrzuO8S+6K4zOOfNh2+28haKgQlsFHe4Y5xr3qdYRxYVv1NBkGLa+/SY1VsWz7fV
X/b60D9pU5lTE5U48lqeA4aJshH3KJB2x6Tj0C4+yjOOW/H4iICiwWZDXuEyF22EuLzME9ebHKYp
aXuvE2y1kMPo+x1smE8ZHp69HC5nRrzPyGCR0fYLOyVJRDpqY7J/H4veybxSaPE+LI0eHHuGRFgD
E1X3w2bKZmvVpcqgLz3lpQKBUb6rzzpPT5gdVK5ysn4ugIvmCRwHl0rYDPdC9zHD5Sc5DsiMORdh
/S6BV4J4E0IWSgs5mzcoIrNqY7eb0xl/8QrKuoefkF3yjbGZw3AS6fgWiyuJdkaWbztyIY81sjte
tpLGWMwXIfrA3g+51junGGz8zDFA7j/AFthVfh+QM+d5cu30sdmmupNzm9uVKUGHwH/8azWttHea
AkK+KAGptWYVZFKOR/8b/9izspi+1bD5xTKd1HAphlaAo5vcI/lM+Uy2iVT1SAf8H77d5Wr/L4er
oN9pY9L0IeJw4PJVw2fyi9P5sb55Rszn+TL7cr+fO2jA+Cokax549byg1F23gWTwW+bZPGFBOfH3
/tY389nAqo28hjlcuREsLD0TzkvQdSqLJc6bJT0Y+6G8r9PmM0vqtovg8O5FdxthhkEKeITq2eul
i21Jg6w19fSTMG1edUGORqGG7Kf4jW+0wMMV1BOArcpDg/h1i+T+ACe782pFKpq16tWT8IwxxuHe
6BntjC272iMqcH5FehwwKAEWrur8Z6LaUR18bXI64PQtZIUXt6ZauQakWr+QmscsV+8J9wUXumuH
LEZW74ldrcxVwVe/lj2Gr3CxSMfXTBUzruzNs0M8fZfQs1i0Jb6+Do3+3AZ4M2TEhrcNkeg/EPyO
mXlGAo/MUaJYZ2EyZnO7ESnlFpuSn1wv5cfZ0sxUV3gj5OK3d/6r2xB8rfyUIneiDdK6oPFZeu/h
iYyrRMVU7lJgsZrvKRouJs9MI91p9Mjs4ZTe+RHUO1nBjjwrit3Kwch8iJxbE3DRDykyQBwOte2j
cyk7c8HAHjppY3/5xnHiAJzEDQ2jT4UoFVGsf1psvwJZhEIgJAOxeoLnE71WTFsPDO6ZUaZs7/qE
2NpnvFN9cLToFDaCCdth6zr37rgQdiaFw2Qic9m9IrPYhp8mpolVtJoX+NMU3hMi76CIl1dR46C2
KjqGNMVtlYBNaTPvdcDJNMdPm34v8OIb58qcGjvTnLQjkx0cVp/KYnX8yq0xPiP5mmJ1bfsq2uj2
5ObYRt6i7M4Z4w5g42NhIMg6AdLSfZaj0rv9HakfGV/8OdCoPcaqhMpWnxJj61UVZbFikuN4fla2
DkJ7uISuF6m46cUo7DplArUMlE4POGp/8i2W6i/FrBRDjrSVsT4+wwF39xyGbi7lIQb37sq+wUB4
3PwhiPhNejTdX9RhdEQPbXlPiy5lpKgbkTnGXSFrnYWZW6oyQ7yqxc5TFq5h916DmphzFIn+WRum
U7IX1rj/Lswu+/AM+olFNb5Wm5jHbK3n8bFljdLUiKsphPU21zG9kMr2bB48HfzbCjWJmNUiWxzG
UBrn98hRPXMdjZXz//iwkTOaT5/NZHONCVsSFghDLyWRvi0dzlFYh/am89ZbcZA+Loti24zZqWa0
7GH2SzR87BTGuN8cznVLw19sUSAAB1KnxErtSS87H05Np1cfIf/IYhsg3IVhR7f/ibC/s0QM1gm/
SkgtbCabN04ifW6LELeIgNmiHeZTeplv0nh0tNADLkmUX2SFoaMK/IgxX9Cbc5Geg3wBuwoP8YMs
pju+rsQmevDixXUVdHMzGCfNBd3iwFzzw/vCAfMQb9JRPb7HQUx6AB7sOQsj2Cmh3iMEv+sAfX1O
MrQkz+0Z0FL9yhN8BQd6Nw88sez1eW0eS8V0pt0Pp91i5FAj8zNOI3TyWipGHAfWwpmArXs7s/n9
oAX8pz1FBAeOVR9h3FmHMRsU/3MLWu92bzTS/3iMqM4SB9xEm7MwPQMn8icZh+ahRmmPAGfaGlKf
YldGDrkZmYtX48d5gUi4oaiTxBKVpU2zrnmZPIAb72mTYsmxmiT1IehIVruCsr/XMIBBqiMTidJT
tD/H++amFP+uzlu9ff0xEIACpkKGCLui8DTbmQMx+UsFxNL3O2fqOD9C2t8NrojMxEwJmPTGB6iC
jq/MniHbDcuGTTgs+usmGxG3CHPvUaV8U5CYiJRA+a2vJOHw2xskrdZW300SYo5SeXPJJSCaRGMg
6q0lyVWvdnhjECRX/Pz889oaO8iHMmymD2qpijYIe0BVA7t1FUnWxgbyreLBY4yc/gHsIRyBMQG5
JT/Xsvx4Eur4WR1dXyQllUWiZsXeUxfkE6OiVrg7QF3gbLQV7IoMRcZWEAwqy1LG7v09l2VDj/KC
xV2IveMbeiVWosG8xchL3shAT3PJ12JRUPdxtDAIlYfCX1/vC6mQZK0r2ZuSxFfPZ4sPdoIlswWy
QVb8N9+ASe6JJo7kYQRvVwEawtL2nncwHNWYn7iPh5nf4zFQhvRAkewf1HFPhzuFy+QZPPJuPGdk
gS+xjBio0R9dHIYJVd1Gf/7anS4EX7qaBN22XjvQr9SR1UlwqjFFch1x4YrxcBxsdFQxOQWi81bl
qM99Xyra8ZCq87ciX2m+RHJq5x7Wfhvyg73kl2jDYRcBznMqc33lyy10vFnJoMQvV9UTo5k0egde
1IZ2qVieonWKiPm9URbyHQz6yAEWCoY3pfwxiCPV/0MOpxow5fky2hgDXo+CjMQgTsfwnZLWcfjw
qSe7BruafbL8EzEq2V6iF3Yi2wbySplcEh0Umh/ccRsoHHvoostGZCkwt5kq9mDr6O1+3OEw5S05
II+/BibvddLq9tQoRE7OH+w5yeoAJOl82L2xYAGUvd9g45+hS4lGbBZqUFuDFYpNpq71exXbq13w
wUTiyQnGxifzJP1kFqhBPPzgraRNRPETsYMmczgqusEK15sCchPnXgLiWY2oUgmI60bHY2JrF2Ml
soa93RfZBDtfX2trctMmlxJkMLSYQclfthlSSSP5L9RzMIfOzG3zVArFx3RBXg7WYcOudy/o7vUy
KQaQB32R25tjrC5w0XS1JoFb72nG0fnHhI6+FhEsFu9Uwyj/KZLtI9OVlPz4/GYpYLMxOqtnAOXd
P3mByGHFptwJKhkojtZ0+AiNYJ3xNKdwOb1mp7KVrWzTH8PpPsAn2S6IHofKB5+n1XcRrCwhIoxD
9wvZPM/DJIIOTFzEjXcn8Qa5EYCNdlgJ3FNtc+eccUDr4lVHmCUKIj8Rnl8F7uvW/EBqlKyFy/2v
srWkzHoztytrPeHP8fgqA6jRNCnsKqgbMkms4F5tgidQsGv9dvmWfhw6/MZBxH5DV2xe13gO4vj9
7jFT0/XYVbf7ATKZx1N/NlK6FxFLP2okBlOW3f+MGCXatxQFchkEljKHOZ3ljW77Kjvd+WS9zxEK
bUpZ+jkOwuPXTCrMjbMoGh4z9svUzZ+V9aF2iOUTsTGtRd1papyVKGm2EGquFiLogVAD92k89kbZ
1Cl0AYmzth06Kqh6JeSVcKuiOSv3K5N2AXxlkeZYKUy8lPAlB3rB2Dtn0b2f+lRiTmrc5QOxf8Ba
gw+dA2wNSPgC8N3MNAllIKoSYcSjVvKzWA7Th2Jz4sG2SkWpESEFn0ugYm68mxgv9AuGgX+XTnCC
0DR6CfbhRqNoQIhFTHyx26cMCEoH+KedVdPFOCEBRWbgGFcmvFsV+Uxc8p1hn/yzliuHmm0JkDhn
XAAm3i1x4ImNDvhURBJ0zb8IXr3IImL9iXgEAaVS01hmgBr3y0eUyod5QRKW/6JMQONVEhYKujk8
iglTSZ09nsTWH8pCHbnUvLUPFxBcI3I32yOsbsytgqSswkXoWv/U/ltJlfkPbx0Qz7Jb2kwPVgPg
Yry6mC/PRV/7Vjt8ACDzi9771Q7Oy+dkfXw02zVaK+hxyeq/K4TalNSDfLbcggh6BtbQTVx+g9YH
jCpPqO5v3sw+raZpWZH9jh/RLeRCdWVAw+Iafa3oq9t4y4t4ttYSgiXboAE+fR+YrzsYoOlFZ9eN
mxLkk6lBRGmjrFdhj13dU1W66k2gJgzq+BJVtZmDJhfO751bxLLWCiMtDv4FIaYlKRVaVXnWSq7d
Vzv8z8S3USwY2GwrERx2CpLFLA1J548kLi4nlYsGiUeYZncT2j2n/5f5wLtYhPiKmgvwyKw9jzl3
f32O32BT8sJWZmhrj3W232SBhyNwuxLoNVSinaQ8+oyQJ4Ceghyfg8z0CDIp4HearnriX1TRsfhS
zXIZuRjuNmGALIr0i6BQ9ZQUB/If+6pLaWf1o8Wz+K1EOQZf8v3JD4gcSOt74mmY0/xUNAuVgTif
+j0jyZG6jUz1merqe75cK/1bebGlXSq54+cNgK75+3hIZJC1yxPkDSKEbt2i9zCBiLMz2N2ThU47
UzKqIUHH+vuWE88PEb8i1tgWxgmmCjz6aYxt6E5cMc4BjoVPlkAsb/E9oz3N9VHMtfDahiblKYd5
xmZdDt8v2Z3AkN3/xqNHQI2swmsrvWNBuLA/qF9h8RB3G2ZGPplwWVauzz81erG5gep9XNlcyKd1
fuviAdL2huTv5S2wBei/eCehDJ7tFpaeBPGyHq0B1gHkJxVVwafdOnFUD+MeXJmv+68Uw/H80JGe
Ec+SshKNm4wHcZTyaSwlkE/2EsMnNdxi4onNSy0oLvdbCOJs3hyqTQBaLseB7kzdR3SZ7hfBHfW0
lTpQEi/ng5BUPuVvD7kGhfR4rp1empOBDxoLyY//yk9aXiV3vAKREU+QtfonSsdpA7dioAU4z/dd
B1EJY4GO07PRBugXwOEDs1lIsHx6BVub/MgrQ+OwgzEkxLNN7KhksOg8IMYfVjL62ZPrrA6sByP9
Aj5NrogzyhUp10NocxZEBkI7LPy235AWOYLnXPWLWmoNun4BF0kLsxtO/rekPnHqCurCKFV6y7K3
LqEhjgNpx9u/cYJ1tbZd0Y6Gm0u9r1sAruTg0GTxNqkQAKyduesnLvM6SCyPaLn17mPIQlpggcck
IgVSXSgtLWQeFN9Rbwf1qXaqfDQ/cRkKg3BJiGhZglD6xZo4hUlibGZVy6wXEQH4an3fquilPCWz
VsP1NTOUKYOX5cb6WQOrxG3MAvEPzq6bx8D+AZYk8QdDckRxxgG+zScHKR3VTTAR0EoOw2N/gvMd
JBRJQ0WoMnRwBgna896j/5R9Kv6qWrXgJFxWkI5Yv68BvMOd74w8v7EfXLKL8rRR7p6djA4oPAmh
H87O1PR9BVK9eA/vzD5uB6uGwF8zEjlhngIUOCp2OLNB4JdDCXDwg5cGt8IhF4iDDGsllLfCqhjp
HdfdUUtNgXgs/Z+cLPuoHe9kiTLo8sUs5HJi95zJfFvsVp7mIche3SOsBGr/pYY4dk+Mbv7QoqUt
V00QJVHOFQxIrvbFXgLCvuiZm4aVtlWFK2mHOTF9W/0wrseqNVvrq6Yls23bep8aBQbDAyM/PwsI
49B3VlGDgfcwYJPNaQFcdoPF6S8M2S9XNkkgu2B7K8nP7Cku0f5MNYn4jBNcPI6cOV1ZWr7z4BSi
qg4JLDBHNaN2xpUC4nzWOAMvcjQ232oQhtX1LXFdJrtW8leIT95AOQOVIQ9F/scNt7qvanZiVW7o
w0NAFbGpXcWAygGDGfxj8UhhcOi0vzRrSKivsCOzG435TK5pSpBxjkFGCz4uU7TdGimT8iVDB+cj
0W852CgA//zASNcVMeGSV1IRcd8k+cnQB6j80SVNTzrzvswvVrGw8KScwEby2qzdT5hQuZzHiU5i
mzBexzkdn3zclH8Necjv9tO4ZzZDRMuTZutHGZsDxOyBRYNIpXEH38IVB08rWJrPrw2hnHUUzE4X
adOtVTkr3SzaGP7N/oC8IG9iAlId5YKTsNxjoehqup5lEBS11Ip7rbD0ozLcLTOuljHQgguv67hj
70nq3joPfaC2hU2KkLnMOGSPWDhBTHaf8A+V4ScfsL/rN1+tbIAgvhjqIxAyUfaPUa5GUNg56BDD
lapBhWZbqD3ACnwYkjZCkU2KCaYDRumlPTSk0Nfzgj7KwdDjEzEaKk1IPSDK9eyYsZ4dDLcMFVs+
zV3GnCPpFq8zX2lgAgMb2CmpZDwRwF035poPwy3oRUHI6Etp4SG/Rj13tcGlbGPfvSHJS+EjoAFi
ZK5swx+cBFnfEzKfU25ISSBb5DzzxDfTYOSwfFWqMc9wSUpMpKHxU7gi5eZJAMUHYTIkUQt/kJMq
jH4VmMc+I/Rp5gtnBlana6ggEV729jHC4rSPcnbbpAy0ZKeAPqD4pB+S6gpCpkXFVVzIn5ISyxbY
Wx/4kyoLUpinCQIZGfppBwreuIu5GuJG5J0j0fb2ndZWswc24yyh7hlHlGB2uUFHWvmuxyvjWH8x
QSbFZuotWfMIDTQSybGob5xm+BDn3T8dnK9W5XHKg0ra0eR9pDgD5J0ygduwtbPYp0C7QDEqSeBa
Emaw5sMxrb22QlhyeBz7YHSg5z/lHR6RRRJvdxXr7dFw8l8kpyad6TOhC9qpJsq2aQ3F5efCBT9N
a8ur4N4Oh4gt+bnhpwGvdTBzOfKnlSmGnK98urX5iCzca4mwE3CwhgyegacwhZQuDjTuab8REjRd
v2G5AtJBMPGyK0P15fjZz7e3ljK45IZgfNGbQdlbk80juA1NbvzDRdXkkSBKoDUT2HHkGizK2ub8
oC/PwMQ0Ma2vxkMivvlLariJyRkWDv4Wxkucwwxg/xPXhD3CCo4EqV31nh23HKM7y0Y7aPOSOUA0
0lQrXcYwJ1SMHRiRLLf7P/NCsuAt+Z0dVDGTg9xtRcyWUEOAjBfSxeSqmk19UXdawwCWB/zTdoWk
4OpKFEapMx6R3TzDOSpljXVgEo3O/uLQL/mHb18GZ8NuYIIUEeECqkcjJKWjYspRLoCoUXaxbX5g
hnmhb3LwmkW0n7HgZu717wjrhBCG/e4HDGNqd+CwVPqsCMD5Q5mLnw3DmX7/lg42OhnMC0RTGVYx
2ByYMqagcxzT2mKGRgrAPlytiV/t8lqlTJVqfk41NAKfdX3AxT1j807z4TItEQgQXNxmpNN3gDUS
ze741aDvnZiJg3U+9Lt77yI16UXhJbhFRo6s0nVXI/x9L9W6OecM09T5rxcLjp5rsLe4EckwbfSd
9qViPz3pwbKIkvNHynOB2CoIGUe2grYCn/oGTM7kZNJrnVgVibcd+sBq3sWvygkAbtkpjg0akUcf
ZvWv6Z4LdVkGOIcG6OH1RYVe+qhj1Yy1gq80ICJFGwDtPROB2mPNhQWsHeWt5SsBNT6tN73FzF47
9Vno0bhDaKqs3GYcsFnBmJIrU6cxfpXIolSkuMAlWD2OgahKG2v214X9KT5dzTYK+JCSjWN1YZOo
sZwS9LMFwr/Psdc7PZfDePBdBu/KialOMeXWan3qNoYL5hJQgvOQ9KSz9hLBjnNe1AWHnNX7ozjO
2/g8Qq1tYw20G8hqwNlZPmoOCz+QIsle8+hMNATktKtJqjy3ZpztqgVVgUzIPtpx7Gnkp79Y6O/a
y4oGtbBjbNEoTDsfgKn+bFj/m7ZrnR7Pl4ujdjhYFpxXKChvxs38Z8Cx3fpm9HlUALZ0WioyWkX2
LOXAVqru0OzERtVINzy7oZzLpOLuwkssNiBYqG4/r6WghHXioAev6mUAKwcsEB5FU3GJjMYj38Go
doBLq5+QFdVJuziDFSMYjIGEU4+26/JShzymwn18wd0C4PHlV/JKECZuFflF0KXXZJHUSB8lQ288
hJOZsHcRmVibjukLoJ4hkJZoM73E/jplgUY9CP1qCW86+aMMg5oGQb7GbqkUt/AadSpsMrVJ5Xrn
gghqdbCDUSbmA5LykCUhx4Pa1jpmN4gA3em+mnjrUsLR7qGkZDCUunMzXsgJUr89BAJVZHqvldsL
6bBmMqoefdO83gj2jQwsf1xL4nx3792JpFZT5bLnjktUVWNRM0pmrOSqItkT9OwO0LLRe8wi5c2T
2LF541JhCfKjBfjH5rgPPNu9Xl6mik6cus/WtXt9nS/A3yv+Ej/GdXFz+9lps7VA9Fw0E9JqKcKR
VR/46PH7ej+dWVJk89zvEoQbvT9VW1mTJz2oqw/5eut9lx4GjNtLICtzUVND+1jwr0lCRXvs6k39
zsVK6szVGPT83Y4eYPfD6lKaxs3WGxtUm7cCZIvqPhPTqbpV4VmHiVQKkEyV5fWCd2o+dr/DOcwP
XPif2kT4sD+K0CK6ZUgxNH/0YefeArskyBBccJ7BmL3Z+On8OJnttcymdD2Vz15oOfgQVxOf8V5e
7AMwnHo5+odJjfC5KRMYllQRmy+RpxiSowNlc28r5BashLEcQ8OlFwaAN5FuBY5w1A6/Y8Pi6c7l
bhnyYnrPXhkMxYaC7y4sCZMuuDXFR4U28glV96xWPyuuids82swG1QBXqxcDbUgKlYaB54nHA6Fl
55eIHDy/PUgxwbUnbnOolW+y0mxn8okwEZbdWO4IztYlU8nlmn+B+B0nlnAgEWAtufDl3M/gREon
+U44yFoPiP9JzjvKOqjUq41dIQATBUmVHyahyCsvnOCpk/VERMaIs+i9cLFHcmEQNre0qYTDZqRo
qomzKQqkyMF2/ByFf7D9HR3UNoF8Zh9PtEdzqkxaRYvAYv5mMTxSO/3tUoGXLXjFHWC9uVdy1rW5
jgmhn6XKCwkt7WkAfu8VjJDkVWTX58KRoL/e5a5F3s01M5ixCSsWZcAABB/kuFvKCNubBuPdtks7
cJ4KTbSURgQtsPELLquKVaSg1hmsivhz5b7xpF+GsH9WPHYr6zZ2doPsRGxXGje4kY40PP7ggHke
rb7DnBx7pq9mbJsWRwCNcwXhocdTMD+1wmVoV5T8I2+wboE5y3CNd4SQ3fDwHU4FjV88RkanID3u
ukXYu+Oz0PbqTrrrtAdm/33UuEzN4fqjIxizAIKvFlJgma0rQ8QOrWSC6wxGf2CO3UkXYS2fz4mh
ghaKXX0xd7aeinC30f0znlHxB/9CTvWDPF6wzznUeKJdg4w7zTYYo8RY+IW/NjbvkR1+/DB2tQUC
+zYhOm2GaewK5bwiTH/8k6JPDBDdRul+FOe+FtpT0xZDU6C2VwuM2Wre0HNzCuqPqu20SDbUiRRD
y7IkGJrP+aqfUhU09iEW9i+v42X9K9cPlwvNWTMA/AyAdwop3qWN8ZWYPSRFS4wv1WzbEfkTtNvf
fOYHjpqgqecDF45t1Obw4W9XyRShAnBuveKqafy4nMq1fQmGyQ7eTJGn2DqnID4LxfOaZRJtQoV2
7VDoypAm4khpNrsMX883oJT7Ambd3ecDIjVTokIM9Lho5AnaZNTOeqFVWbUfKpUSsKviBv4Pezw/
N8Bg6AqNh1mCVfxQvaFe3h5GInFoA6Z0HOTDov9AcA+kCa5EeLq+idkYofKka+fWNoKakEKuFGrm
Gq4wlxA61+qyLcEbyNrw8ep0guEFuA3ycwDxRJc+XVAmoGToRtBHf9ozQmDCNyXhlrsqhoN/fPmi
/Wbm6KAV3PFg2DWtKke6Knr/xaSzSePEgNuR25pHTuOxSpoGCsfE1ic6kCN7HkhMcOpfX/4X82oO
swBwHciFluFqIzMfqqqLbOCfOAwDKY+KH1AUrAN5kTBVAnHmpMsyuwAcO459qeokRNz5Hs8+Up7R
LHgPnLUgC3IdbZTfyqcmM97FW5Z2M9NsWy8RqBxiQE6V9LzxnI5HnDCBec0uku3LhWPMr1dbCtmb
Yn0h4wvqGtWAarVmseb3oewh2dYrKn+y4cshYuBCqKytcIKtLNmsYd93TGJkRCkRZa5J+3XdHcZC
S39o4b1N/+h8eHrbz/8gaT2cVq+Bx62gGlt2tzcrFFEC7k4AIjSF02cJHKJbQDsZgbSGpDrQ2O5H
g6/tpRmYsxOb3ESZUSyMRVP1jpFbndzPI0lubAPCuGMmXTxknBN/C4ljTNhyOJd/dxF/WkEsw1Jj
StkDW1T4KE8XSaXNA6L6gUyowG7wGLuuedDsQovxQP684wlk8RdqhaRrM1Nrm4himsvXiULkISVB
cC8HS82xl6BSK2dHdpKrtivfXbOUk58iW7sL1hwUYUzf/nobqTB8u0uCmKpE8FVqALO1nod9mfMp
54sUCWLFuNVdpNLqWi+kS6lJCPeXepWSjHcuvbZfT+V4fjw+xGCp8YMMID1/p5NDb12kQJ2MD4rm
FvfxA3SlLk/T1qzyf68JnNxZYW2eaX88+Pq0SjNKgfgASDl4qJqpy2vU3PKYXSS+cLjd31lxgl+i
RqM3WNXkXcISFtaf7fO/bEUok/Xs6intCC4fIXlc4RhqnVhjYwPvyK0BG13iTktn0RqMOSuzoASS
/a7NYswzK0kToaXKQ3vcqYQ0nRBvXonoI/KRgG52hQx+lhNKrDsTG4lcc1KcZu4z14Uu5Lm4bnm1
jVV380rwsJrATeT0mtuSvyM/zrohSU6wF7vCTybocOcb7HeJvXuL3asoLMpxxYqKiFg5K4Z/nYjM
hhcAkUFcxgEOMSxBuXtZiux/jepXv42ZhPuHDGnFNCBqb31HNCmLiWszyfN1WjFx3p0ZQgwotfgf
+uHAnaFGI4cbgFEfGu/LVYmo9zdlxDTPeZT0woQCbK/DAXDDwHT/8ccLSdfPdMFRQwPybTrOuOpv
AaVVYBQbtqwj/kI5sZeYM1plGNmNhVACHzEig1MWmRnqjMUeltETl2o9rBd9ivra1QE2sx74LbgO
G5N3Ev8tAcBbyc3pWH+O013WWgFcphQRxgHt0OqFU1+F7WJo5eYyYqMKgQ48osZU33lx+y7wRnSL
o7RJi7Tc3KQny/XKP8IdVEJmCE6iorm39d8YO4rkFW+RmFiaJ3f/0W0d49V0klcJ2gr6LJ9j7Rq2
K505dr8K3YpSJrSWTrdSME3JpWM41GSslqPSaabLRbE65sv8izLI/h8e6jiaZLYdbta66eo5oVPS
4b7g7uGn6IskL+lSGUf0Fh+xolwNpBaocBtyeCz6AoWxN2hTvsvF39rqaFpZcbPgXPe47AWYniT+
lRoEHZz9bIFjyrFzClKE2tQ1jXODtCGJV5VKQ0d8ssyec+HwJJ49Rjku2KY3mQmuiplcJT9QuXI9
QBRFZSOCtxo4tc29+zOMyLf+A28TUlfp875tSScFVNDM+fTG4Z/BA0EtNQIODB6PjL2xaRwU2J2p
toHLqN3Qt+QsIVEScDUPpyAk70MyVyxwud52WMWUbpynOFXdCAku0aNn7cCeyG63/dJKbyM0b+rd
aYPtFwTahM/LpVGFyqEmnw+6lF6KsdE0PbRcIXVk0EGfkz+73hcihm9pJEZ6v1EYXrV3XNVz8Y0s
c8WcTSqmEdMWiJnFnx22Ed/+6EGyMeAf/DdZT5AX+E96GyhaWwIxzwLijX7TNKrZbQJVprxQxqVP
Wm26VXipH4NXL0ysTT2Xn9ngwNUd5eJ8QvRJXwp2av84w3bIJjE2eAyaVAOGchOmoo6hF3suKQN4
u1dJVrrSCA+2gSgOF0kwtu3WqKVPtGFLY78kOK8E6KQvy4H4N6vSrAeIK+g5Lm04paX78apEISnW
c2x8DzNC3mHv6/FEjE8A1pE01mqMZk8rK+mV8eIlCZF/vgzb2565aQwObeksGMAT6gyo+Q52WHwj
f/p5p3jYqTJ88LkordPhK/236x/FvdXOux9jUEZ/WTpxoz2tLF5yMqKTdUv+YhyY8eT2dZSgaHGE
fRiyMJSmlXhoRDEz5CrzflzgFSNzSPLl+68F22q2dz0utS43akNZ1MlFqVcggDKXSflYzrMadeti
FqN+xi985LfOugVkRzKoEv0r08YixsBySW8zn42AwRBUZlCkROWGQkPvXbVtaGGfhqUb6xG3ehBR
49Bog+HTdRRhiIElX8jAGIhgkxmXsi81+CJiCFRSDbZR04i/PoOxiFaxhJrD31kBe6f8pzqy7651
t8nXNQ2rSk0cvhlH4jr8kNYs7uIqypkIWvYGFsJ+jujiHPd8Dw5BC/TufOxZSJukgKO12HQnZpZo
ePRKIRmKKVXZY3BSViuIXUylLsMZFUd2mtJ9WBqfJsEkqxwQSOBqCmay8XiCvThieo0wBn7bVafq
MWOvVeKpsLFQZqNNE0X6+GjOxK75U0Aw9lW462ov9Bc+3XrmF3z4dwDYHr04PW+aJ5YUeb32Vz25
asl/kymRmwLtPD5ZAg5O+/vHfup2BlrC6F3RWJBHZh8sTJt7mmf6oGWMcd4i2yoWeMqMxpLtpwTU
NcWGsUFZ2oXo3/1MlncLBVBvoBeiiQo5hr4G3UfuGWUzYv5bBURqvnIZaOYXj0UMQT7lbiRP70C8
aGVYSC/BW2WSvOZfN7yNOpaBQl8Mf+Eu2890zuR3/9Z9ikkP9syawAPI6R7Bu9QJTyOsZepXc9xw
2SSJCOb84kga4vFeCSrLyxMdKFRWyDp8M4sTIHpzl7rTlIOtuN0x4EZqoAnpMhSvapIICulxSLpX
O8wc6t9uz5napGoDW8VnJAcD0U8JNaFfHQTz6WfllUhxk+ZBYpJQLqTmvYUybBBG3JnFjjJxbniK
Ws9uY6lri81uoiP+hq8HzLm5qINO/H1dt6SuzQgbPTpSqKgPcR5AWxdO2g9T5YeSeocV5LP3JBNx
51ezDVGBum/4197G7G+1sT+I7DVZicKLKO2SVmfjbAxqSkL3Epj/yyeYXs0VoPQGs3ScXCpbtFqd
Jp2t/4Bo6+++rir5GD3+QsGt+hSzehce3xRRBHuGcXDIbKDmnmJ0AlzbA5OXxWVNuEA33fCU6310
9gY57jbORbOiELASyhMz46x8yEQe42DAwAy7GklJfo7lbuNV+CpaCeA09r8O0BunZ4LoZXsAEKIB
emiRd1SWlKkXY7SxPghYpbkfsrL7VOa0v2ueKgNq0BqtxK4tLCUm9kZtlQNjNT+qrb9DedLKwHpT
HLG542qx199TteKEOBNY0p+HF/MMFAqwGV4cNaKJhbds/8RiLP3qzkSeKTA0VDFZ1Al0xAdPG1cA
AHyqqXngnTmgOYf7k24ue6k1jf34Jstr7Fani/Y/5suexhH/3CRrWMxOdc5EXDF+jFDoKKo/ui8J
sy8Ex4cOyHAc3tI95lVD+r92RJy3zsTLno3Kltydwa0PtdvYqxmg/8xH7njCTyXyEqht1qM660sV
ET8owCmUhRe+f14PzXTFXyi2rCVYa9D8y10yrFSHBsuBjF0fyoJs6j3rIo+NV+cz/5i9hTPIBoRU
GnoJFZMvTvGfATXgvaUs3vr3rt4za8qeRvfs2PY0i9TaBmYyQIfd2FnhJBzTPF0Y0XpqF8WEvHo2
diqykW3Edhm/GOl5MgcAqsxdLSY0FQAA8X6m5chzKBwEKJPtASWz6vdMkPdWlDHtyutdT9U9oLSO
eYFcMv3xbwTIUWw3+gYHroZD6yRcp66p7Y04UON+CgMZtyGy89YkmQYzCqgW4mQXFW6j0Gy7f5uQ
8Wfcnd+kBKegTAho9oWMS6rePfrISNGiA1Kl/2uXM5BIvYYCT5ZsWVJhClNL8f1zbkzPWnrvgWg+
b5yoegsb2JaHAwmlF45CtoZElJ+dc7TXrk+6WqfWXBPGvSNrq8pz2CyNfSt5ZxiC6fF85CWyX+Fi
Cxspg1h9wwmrJLDotAqMWf4sk9BU1hWUq26r5foBCNTgPkNH+PpCYYgq1ZtZyMcRDXi9ltlKqW9w
DE0MNjEvePFuHO65H7h/GQql07Z+0EmvW2ZtiSGZsj/Xy3X6q3feZTOQcU+HeBmZoUuJ1hhmX0dE
WHs1dU4wGkJRDVDNXxxv7ZFPrsWcOJAF++P8HiKUeZTFWuEZKkqnfOaZjLUHUCVNmNOE0nJ2tBRB
pafsdnFQxEZkNqaafaMChi9iNdumDDUc+RFsf9WFqhhGMWPEkhYj/l+yrCXlusmxk0WDK2iL1c4q
CFkOiiniM5v1TieViklJUDqwguILfakJrIS4zH0+vbz7bh/8p52TbMSJeLn8CYMw9nGDyY1uLtYU
kS+0oqjTevScfC3vvaFi2CfCtVJxYqLBqb417L7V/IEfBWBUCeSVc8iLG+1sEgWdmYrJacwonFVO
UaOM9aWncB9taoqtDVgAA10hPsjg5pL0g7a1Ypm8mYSb6gkMsHqq6TFQr3Dvw7WGvThDwb1HyhbN
xtVBgpw1B0WwPq8XDdWEv6RKTtS0xZq39RmStHF8oWAWDLGbW/ogTUhLqFqEKQztNQNEQzDEJQKP
m8zYfKThRRcwIYMF3qT96YzrQ8vMjjP0UUWDGmvXQBHuDQ/6kOHM+53VkEiedTssRHZpSaBB4UcB
MwoRI0DXYvef5rhC45DncFCUj0Cin/tNTUeeQIV1etuj0XAz7C/lyWxf4u/3D3xWcrpe515jgvoa
Nq/e1f1xnmbJUMYVbKM0OKmHUBHu2Fb3coK826q2m4cuVSdPTNKoo+LmxLIZWn0DJs5po2fPwU7s
hhSSDxCg5EKAMo2a810ogOOGFPcuThbNJJr0TsZzDARz2qZwViWvPqeQGk6DjuDE6mmr0w9uI5iO
vsGdcfX78lXGYnb/Ok5gFNKCR/sBvs67e63kXi9hZ7o0cXcQCMa7u7gYHMwc4E729fWkLCDGjphG
rtxRXPqEdlxSbl/SMgVWNVFyw2+oKNcoVzi+drOQkd53/5xKLStXt0giEww03jiN+fdx21OvC4+e
vIhQcR9dyKnGgc5PAFAS9xUBdEx4ad0ZI9Pdxp30mfrrUJCB1A1VyR+CSOlw/iQCs73ckhqOZIB5
irhR+T/ECoswbMQO8S8vwv9y5MT7KadB2Z+1qMeo6GJHmTa0YivJ92RjArtCbAJ7rBgOBAd2jVgy
O+GfHs9kyPKrGNtXzPjJTvAdoF2R9/4wMbiCADdSeK3BEhFF6AxUS/us9+k8ifO9PAMHatK6rDTp
cN9ymtBhMyXpzhrCAy3NkocHjeydwRgvxniDMH7GyupR9G3KD2A5hc6OH4abi35bTJ/dHYWrqRxZ
JoZKx/Ubnzxq1oFMH+NRjvZRbhwPv2FXkGV2rtovYC3S4SAT4XLQXoh2ckB9xJuc/2st1IFOyk8p
rRFiWYnRsu0t7oYpViro88wXc2JjPRmy/2W/eZVa5PzUZc4pL2zyLZoqRQYgbmjy+FBKGm/ob1a3
g026wQ0dTMl6Y+OZPgbAFB3gns5CsWqH3tuNshblUjSohKnN46f8SXWK/+ioXR+O42+T5Wu8AIVg
u450vAA/8SAxo5R0D5V13jPYyczJJcwiz1hzRdAIRscItN3FBzqxNutzxgUxswLem11zE6v+QSfd
Miqp6c2lxH5XgCMZ8+JDe1GJz3AEB1DlbXEPveo8S/RhDaNm4tgdyk+ELoDryQGiSS/wAwXdZl2D
CtZGbePC2jTsllu7Lf3vhOCpQxZaSiMrWK8aJklfAx23l54SYkRq0es1Y6QAUVM7ehtJAlZxElOO
PFT98dqFc7fMXnekSqZFfpUjSrroKePZkrqxHJcLK+xEkH89rLeIXKA8rGxKPQRHmDH2mdoZyuQf
RGnJicqeHrDDsMCNaL1ei+EDQMSXp3tIryt/jEHfg/zAMu0oTwlC5WcGzH9ONo+HNeUZpHskmmdL
TzoS28DP4/rJQFceOthSzYKWe3aKs3lHCfGv65qyw0goxyaxGqGU4Z5BJ+8Ow9LM0dam8IUPIvRw
JxaD59wFCreo1kzFMVN7N368sk2c1BlmINSjaWDq18+FU3Ptk7g/FhWVBrxygVfLxqC4szC2J/4R
3blsAW5MgErUGrtwVLgegVOeEHyTQsIFiub0L1gSnDOvZkuojnIXmg1Zk3n7RE2FQ8xEMi6jEOAV
BCkFrRvAK2323mnNqirMBdQoUTR/RbQX+uHTrrqmpg2UWP6s4X4HqIE+HsonBLYfhLDrLuAKnims
4vKbq/5OZ7HAkipRGM1lA9pMHW5/7I0QrVkn3tsPT67qmeF5DdKjRBfrhRB72BQ86oTb92Eqp007
RCIfqQKTI5juMawGyiV/ME5osg6vvL2/66bnBSlOggle0ic+bgRJ9HOm44y1ANnELQLJQv0PRBTt
8Se4koYoMQ3U2LfrgTUM4ISVR5XfPJ9Bvsyt0j0aDdim7M1WkP7AATaJyz2M0hqGvcN3Fqdt/y+d
UEtGt30hyk5WazuCsQEU2KHzGCXTLmAEX6OTpPVZpjkI3M7eTGz6Krnexls81Dm7elLXpX/bD+zp
0SEcQvd0nyOKdy8qCpkNk7u0gNY3AnMtDmSFfNPHDKBCUqqn4P/YPnOvKoAFJ22pyZxq1AUxBrFs
aL+mOLcI3Hed90V33ixG5pRzSOXM346JUBm9B+xoO/bxTk6RfkPAvT+xpdinqcE+u0DiYXxH00EQ
mEgyfW+rPDwiQ7vxO65+453NVYkz/XWdu8tYdOo2QGhNbdCRpNIh1fptruFDjBTwuIybZQiyBSR8
vA4lyzYI7VeF8YiT72Wn3gh/jvv3zJ9kpxy0HbVmOZGx+olgeWzfFtlELPPLFUcAxTQvGr/Quske
/Q6sCnPeajfk3xXtwTWFIsMYiWum2F7QJZzCLwgBQvKZjoHsZlJ24kOkFpYdYCLYHyDjscv6ok4M
PsplPfLPMYSZHIpTneOsp1rO/pfXsihelVejrjQiEG+nnEl4/5T4WHtwH1xyk0e4nu+fnf5Zq12l
tdeRa/IcHGFw6iZSbWscJdwuqHn5pIUiBgXiT5/calrLhrFO7vuJl9f0NlyDAvrWjAeDwy+qtcAH
FOn1aJCdYBDg6jItdR2Rsy+3Xd59rrKm5yHK6LZQyPw3ya1pnOcqvkAgXLJdSEH5tphDHZi3jPbu
/76i735wzlJCiE6C2wytCib9Fa9mWbL1YhFyl41mIL+BRDUZ5jKa882BH4TI8U/kHs8CjMmoVu0j
4aIJzMZo28NQU91O4z8qUK3i9D/IILVjJzMHNGp02Yr59VtFeDMbgVfB+5QBkO1oq7fDDUeqIkeO
0ey0gGGNqlEqAP583/bDFgq1SOqlbCCR3AeGF8zBnQ55gvvH+GdhPIIcOPVk/SMJh2cnCMUdIZ3i
NJzrJT/l93aJT8CI3szBKHiJfrGIjon1hfbC5aczb9VeocVjgUgfj4u1dximWAGIcWpYNSHYh6Ls
mXlCDcpErQ+ZeHyIkzGNSLiB+hHaPscAeFskwptyZo33eqD+kTJkxp7CxcTKCSV65mgQucuEK6z1
i+tMcXyO5dcsTp++ErIJA3QvTP3J41F1MwjJtrFRUGSUVKKz8uq/OSxuo2K8j18Aw6Kh2nZ41Urm
KQgrNG1lfD4cU/vJPzNqr2DTCJu1TjAgZSwwZG49vGzYqEeR9tvQzhRTwh9xbACFBCBdsH9cMXWj
Gu7nJ+d9oLm9D0uKjelx997NsjclwCaCgyjCC5Vz1VAwib5ZJYx+BKTeu964YXaZgkuBG0yC38Ou
YFrzYbqSKVYrVRzgnhbU2QXCcF0PKLWwxOEoi8cUzy52m29kGrFsrQBWuM+sYNwGD2evfc4viKZO
7MibYKHdIr3B04I3eLxWIsHQYZ/ZITsMy5lStygQpEbqK8IlHCViKqfBDCHw4j7/2rewBfRSueWC
goP6iEj0FceRNer28v1HdpKmSlbeyS7Ey08CFaL+Bwtc5Sfo8clil6RuJNQfBQTu6IVcj906YnQA
MibkhyjmJazqVzAz3yAbJUUj/TM2G0LRgXTKWHtXe5KglqTdLInGVKy9TnGmIvW5t8zMub/wKaWf
+kPoaz6pUteCyWth4HvYO3aMHGSlk25Q3+hLbkXN0MJTV325IA+0qqw0xUSrNIgg0jrZafuU9DKl
adSA6K8a/jWVUJyffB9o/vLnpKbgIJQS8xqB57T/F+Rqz8BZSN33SH9S3Se8yrq5Ogi0p92FLV87
+uicOJAW/9xxn9QXOErJtK/rIq2QHE7OuEp/Y33HmTabpqtJtt/Is0a+bfSjeSEoJgs74BWcjxOo
lGf0EyU9rIna6o4EN5YxEHxaEEBblSymFzuGGn9gccdfYqSZ4R89852OAcghl6lO3XmNJy8fqZ2f
e/os10jil3jhZ6O7RwVMjbweo8Pq/xSZWS0PWBzVh9g54vwEwlFtVhkHag1flTYVefsBqOXXZmyp
/gjETDhLDeHK3rG4xn/kxCHpBePSQ0VMSWrOycR1aS+bZrMmJfrWivO5QoYQc3+ZqrPDuGO2uZzV
MQqXnhVlgfWE80ahVDFSrz8u6xb3HqDXqdGiXa4WOskTjYvMiMbUZctwcZFZKd4e1f6SHhVjfHil
ytHo7pnous+aSSEnFDo8SfLMdyCMgt5xnBWpf2qxNneWFStQ6KB1ritV3TTBliJFnqrDEN+5bcH2
tJdudz96vHnm3/YyvisZdZRng0+7XpMrpfqraXgnF1048TiK6B2wnnJt1sLxHBUt94Rhou2Cx4AR
6mjlVN5sNlmfIXllcaSiX42iKoucZjdZ92KboHFFnIbBB7zxPyIRkvu2wYsJ0QsgqueN9iq3RzZo
CXdnl9gsFOZB9ToRWmpsyRK9MCWRTsMYTSoymWsl3ENPkEAjor8aIm+5NPKbJzCuB6R8WkkjE28T
u+oAwZvVeoxgQxIC2wB0VB6hBygClLTr7J2cEpcMdDcorb3g7mA2e998HZTOwHNc0+kyiaWnwzkQ
liGhL6lV98LPkeUAgQTnfsRIiGsF6sCt4QIT+KAr6IwwhR28ri/PW67JQiUg1Kr39poaZqO63pJs
1lAXOSpfJDEgU7DWkygsRUqvn++E4CiPhDDSjS13lhEeI+B6Pi7hz5RVNh9F2mjoNFijAZO73YbA
UsAw24zxMCKcF6uKVMIRZEoqPqE1WEIYsFJccer8yAnwJhh5Ld/ulx2Rr9OGuPB8kW8zj5fOxuI/
BEVpnxbI3a4rx0c7CGoZ+1azG5+e73SkSdOX15vIdYJCoaije3T2G1uT+b0E7ZM4/4yEIF+WELlu
njIRk+GVG4Kq1BmpvJIOkN4HKvxnL94oDXuXKLirOPIIRhxUQ4YX+qJequnB71TtuRfD89MaBHQN
8d6qZ74erPMVwhT5BB1e+2LquqGy15kDIn5eqQovsBuNDlRF7TWebKIOP7fH+VJCnqtRkvT6/v9G
4xuXfqVmsGd7+iHW09ePwqJZA3Num9X51PF1IxRhrRIINuvsyDKnd5pg2pffepdJlfcTJwABKLcx
yycsA5qhhynfIM0JmcAFpnu1YX8QfKtn3Jy4Y0GT5Q+ZvyPOBpPPIaVn0ILVl8bfoTI8GXYuSY3v
WbgNWet3QZFG54HyeztAkCldnNQ+7W54fx93w+7DGrSqrTcBlXKS6EwT7xkIrKN2GOZzI+WbsZ+L
ufyZSlJHkWaMQPak1+7y4Yxkp/4p5aIelpvREYZL4KlEUqs03X29ybS24/jT460M/yJh4yunTCNG
BpHPiU4ScLS7yXRVmwPHMyBBLz3ohzk+fRGcEan1DfK6e7FY0qJ8WP2svjkZZGbxsfTrX66Ysbw9
mhDklXG9wIJfK7MtcmrrCWteZRKTCQL3RuWzLpzYU2RXeop8LPmIhSyfEDisNEqrSNDr5V+1CZQF
BF1dbXwmhVrmydBNw5by4PEryyvUAwVFWj7pwcPuoeSbR13Pgi6QjUs8MMS+/PlHw4zEvJFCxJk7
PJ3MnBJKF9aOT7oBmHqdZ5qt0j8kzEoncRdysa9/qTZkhCpYLsZU5fKw9qkigVcLv9nJs7Lh8FUk
8wTiuQ8aQWGODlM1dGDEWSxREh/8GcZ2SkSCERZd/ahX7WqKFA2Zff1Ise+2mT/rMGeoaX9ZKDt7
wiYyjhUiGdZxvIyPfMi/cRYGOyrZdVHavPH3brSsDmHqPSmJJ/Y6keK7fSh1JVY85Ul/02qCJz4O
IdrEPNA6ePRMzFCYHJ3IWyPWFL8DaA3/WPpePCZXXwiSdKwxrJ9jm5pIXlSM3Fmucn1aPqu7QGEX
9soB/GzfXFN/MprbUODb04ERy4We4acXPyzLZgEL/0fjJt9+ENfLEFgwHdMi0dClWlDVNKwMNWSi
2yYRsaMlVbpqWVnOhH3HkyaCJA2heWKB2IoF3CE9bxM94kfju1Rj5azmwDyg4bPkX76JEsnvYku6
QeTkdg+igjfu1x+RwB0nRJUCTDTLEnaRK/hKkpVicqXtZhrtRA5x6v6OohM0g3c6bdCopyGhLG0t
WPlLY23l/0nLJXiC6i6XOt0UctNJQpGpgKf+6RE9PbCqGhDea3SdDak7TAmvWhVeBotR0mDaJVDt
JhDn6JBTOmgeJd662THCXFzueoM/SsWu2AXiWW6rw7KqQDbBBSct4KACUvMblYM5YBNJY1Z/SyMN
NLi4oLqRnDGrSdGFjUoZ4qQse16L0nYb88aMV/E/3AHy8qpsSVRJLDJGcTVRQ7PST59iveNpuK5U
/S1msNKT5mId32c28Krc6dZrWsJrI0eg+wmeE8xtaCMq3bB481rlAsRYr/aUnUMfkL+aookEbWJE
n77FONfkI+XKz7kLWzvzoxUYEjMVvDGIa5pE+18YYQCQvdNC28FRw4noWiGt2YsioMZoXfhO6BjS
b2ttXUSw+41hJcGr5nHRcSvvlN+oleOrRYDRn3uYKh/GAUDO77jGExNpIrI+qeEDyBUebbYuWg9J
X7/He7tfL/J/136UuKjOGE0p3Yy5q1SkvL2n2BOohAq16GAU5v6UwY3YWOTIxHk5nclToknlsRE8
9oPwhYbJRAV/2MArdPP4gawdevIQ4I/QQwMjlHCGZqnUSXYLJDm7IBnpZl61ZX6cX22tHvPHp8BK
vmruZli0eMoV6UORKo9jgHQs1v7eOY0w1f57Ux58TcXNiUDyzvVv35UTnDFLtOyPWh2/HQ2Y6oi6
j+qa+O6zl7tEghSNOTMzYhELHx/TnurVK19SQAUvBrXnEMzejJPtesW5f4EfrrZoR8310js363Ms
7ViFcSLISxNf4lzfYYuvZm4p12+7h/zHWxQ1i6Bn4Zsans9jCw+kKWkdepRtj/qZ1tbdXXuYIjrS
xXwo6NXDY2yU7X2xaCfoNuN9uEPlQidhqowSEpb3y9J+GMtEylddq19XAc6Lqii51wK0nF356D3P
fQjA7sjFWB3eSbIioh2Rre7G5WSqmAxlM5WDq+A2VZoSnye9zWzK/L6a2X59VNiGzzUdjbodYNF6
vyhsmfphLij+FknQNzzfkQQFA+o1vKguDb61yOPIGS701D/gFsi1v+iPf+pmq+NGEUxEO3LyaZWm
iMZxh8JiC3jnKz/3MJ2sxnEWNN5hasAiucHcp5nuAYDedDbSfYrkFMfsi0Asq5njLqrcFhIfjz+h
qnsZc+SpJ2BL6w81ugLdjRU1X69Ci6kVcehwOKlmosGXU9eBCp5HLzJ4EtHDw4RtAqLGPqBlIGNi
jVcMBi8wp8/mptjNXPQ9mXOfZQaQWbVF+h3mU3s+FwQ/Ol2LQFkFqqyy5CprXFVsxAAOuLypiSS6
pZu4QsI8CRkZbX0srS84qyefOWHTNVdwHp7paLo73QAiDYOzYvgm6a4kBBsPmZhPemkyPKELuRro
75RHvLibGDBvarEgKdUWqqoYJJYQzVb7SjWeEh7SAafpwYlKNWMMcxmWKaypeZGRps/MqJ0uj4+3
R26TVYB4OTscAnJ6iy0l2UGiQZnTS/quN3rStYdJpCaPwYXY9kDoDPLfm8/sFNc7MgNFZ5ISuknk
qenK2K0G/6OQyK/XfGIzOeObT5X5x4Utijll8M0NgoY0/IvJWYGXZ2RFKlfOx/AXkUKGaM60tGgi
eoDSCT1V5SOsXClB6lZJM7lgbGyP85VBPAmvoUdHoqBSAgKVpbu1YNfR7/vY1dgSemGC7NgI5OqN
r13S4Rl+hf9htawRYQbS3SejzqIkPx1t2xG8Pv9NiT2fTeH6hPRKka3w3tI57vhTyIMgX6iMt3fz
bRrQsdbY376FDv1GyfwvaQdHU+EUPwjyLyBnzUXrOOh0SJs+K3zMs9qJXUWXBnrRXdm2u1gc3Ugg
bnQhc0G/tslGgZH/vtlAysvktLnIGcmL0uyO3Pdu9A5tv+tVR9o7zuZFLpn5Oit+XFoV6A0drTSQ
IFv47K75viMWYmTd/wos9ON0LLAabdn68cq67HAR/B0H/GL3x+PXbfl2Yxmbh5jZ2JrxTrT2fG5b
Cp6hJ+Q8PUDaIMu386K8KuipIjwVWILrQGDMFnPuLW45NvfM7jvz6TIDrmVi6D+TQcbwmyE+hrUZ
qtAtdNPzurcBj4VMNpUE6hOlrC0jk+jbpdcZbZVXZl84qwUpJB1b7rDi699Mc45GifvCTxdZqmXI
8Q34SMer2nKHOS7jamofBPa4aMgef2Uyso9tq/6XkxmsD7PvYIhcnzBUtJtxASYJG5CNs3HaAh9a
595Cv8htgTh3FVvrbiw7OzA762CGQdhiREYxseQTSKGtkhkYmD/fUPNSvxZY6Riayq7zsknTyXaM
ghXvl4mpXOD7N0SvPFB7BGsgSSBFFPaO9yv+56DZVQr/z4F7WazxJEVcKs35Q62fZrSyX+z0mW71
dU6pITo04ks7VuivH24U4ygJPHUS6+OpqkImcrplPGG9XvawuiLQmk40tqQJIWs/qeOolzj5mwYL
jC3hKILg7TWZEJkVnZqfftx2ldIit1j6D4OUNXqEWbqL/XAjVUDZgMsdi0hzYnFHruESUbERI4GH
o9DCG5S7ds05wkFXKZ/7gs5h3nQsjMFJM7L1IMCht2/wkZB+j9GWACSmC5APt46iSMCmW57U05kD
I/jjagUyFKaxj9a1kzNl58EGbP/ahKdOcgU/69LRk7b94dE0wo7HTjwGgsiXZ8z870afyIIf/H/W
X92QHElF8EjkKsOWQ/V2tAqm4bba5grB4J2tyvL6AGQGvOiFOAoH/pdbRXa4+u9Fg1Kkh5PSvcr3
S6RmvFI2e5z0BhvIACEkHlv7DRLxzEBsEXNalBaG1g+oUAOHurwIwPK8mHYjOQrZfSn6QYlsHhXO
p8BY698AwLhizGq7jwzmCotvD3UnsVwtiRpPottT8MWCH0kyhKsarq8B0aqEKdplsPiT05hqXHnH
oihnXiBGHTFHZqsrlG1LZ9ECUDTwr+9pgT1E5l5M/6unzEehqzU4+fvDBeM4k26NAqu6/VdxXc7D
kt3snF8YkRmwNduY4ZNLQXF3uRDQ6LxYrxxReSa3u4yxilo0cGQAwH5fsEt9RCyurdkmphh+UTEv
qK4fPCNGxe3tsHr2RdXYb3WUlBoudSHzzQlvc+WguaMPRoZNoRfVqytm9hdFVYKiY2B13K+0T/XD
Er6MSgW4NZwvt9e9I29uA6zqkJheznxAAr6yizX/nYbYaKFb3aTlUpyjBUrRwwKWJLB4iWHl6g0H
F9Ho8f2pIVABWqq9pqqoyYgEcMt5IKTDOxmsA13hZE6AVKfFN+XEzwsQqKwuQbKHjZk+k6V3y5bB
XfST8aaQxCGlMDAkLMrqvX8w+HFiiWipQI/mF67IG9xuRi+iY8wDUV6iC5ukXAgf/LlyHDVnvciJ
9AkejzLbO/gUqJ3LOfeK6aj5X40YhKs17sBtAm9GZxLHUWPRrI4enW+pyoeArM4uSJsChMqSHC4a
1C11wkc7U7UZca4Pimft1j29yGSbdG11F+lj9JHpIhRrXtqBJl1PVPTVUwEI8PVFnaFnsEAwfuUs
b+Lgc0Cc/z1/LiD0etYbHQ8sozIdFnBYYw9X231utxrRvarI9nL8m+r/aD2k38+DMWyZNVdtDj3s
Li708TNsiNigHRMCzXXlqyyri1tygyCCrJPsUbIOHAA8OrFj70/gIH4BQp4B7KHyXn2Q8CQqpIP/
4LpUEhiIwMF20+/qaEpf8U4KDx0LFqdniiJo3q0qKdsXZ2+IH0uY+b6ks3+63uCM6zMPWYJY6BI+
FQhjZbujofToP9/77ApVNCFrf9ffzZkHlrulhnYS6iH7wFq8KYWT90ETHY+N2uUAHOcSBhjeXo3B
EGeOGMTMCAktetc9i9edfx8xpULiGaFEb4WCjE96rIpy1YNJsbMyHg0r18WeNtiZTzWsXZefM/6A
nG4FOc2xryOdmFjoshokuXVmbNAR1yiqXXV8S6i3RuQZX3IiyOfToE437bxhp+yK1H3Oi6E7AGbX
GemP2+7p9D8RlTUDiw4vPV4uugkj6xUwtorLw8C7aDVKa3Y0bvrnmoTQEU/sKGCWhGkhrgJmxkEb
6QKoI4vYtUyATUN7TmK4qciuiYVEJuqZ8az4qwtZdUft13tYRjAGbhggD6cukKQveC7LsFOF/YD2
s9UXrVIy6CDr4ET2FAEx5kKW4DmEigcCshUd6+u+e1gRObVQOMAs9Jhxwpia9xcNgqwQAMbe4iSY
mRCW5j3OkQDh4KicpHuop2un8PC523qqFPtjIDRrteaQrBauUrNI2u8F/79hEQ+Qe7Xf+SC/tHuY
4apugH1Ld2b/Nhc055tLe/nzs9OJdZQmhPGgdrR4s+5X3qaS2clPpoueQ1BZRJzCjKEHr7SpCufe
+t7wx+5+0jutDqmjuVny4kGN0Y3yD1n8bq5LtUMlVdyQS6TclpATOl9iJmwddPwWtjZxBs2FzbFb
Bvn0CmMEmjFqlmX6aZtnKP12G0c4UOj6PsRdf8Fe0Ky0fs/wwD1FCQNmEYe5mZu2mbaGTezSmQKs
RLMnbJL3eQ+YMsFd6IDfQy1jMlH/iRlne8tNJaSPeADkrwC2QeqLSNPxqWt2JRu4XHEfx5CI3COX
mi9+MlZY4WzOJiEV+lWxHf2BXLnu2F25u//iTMoSljROhkVK1Ia6dVYZolwaHxCA2iYmuxh6UQAx
hvvRDAhCwQNRz3WR03kyEpK/A2eUdxugOj/BLH4XOLVgeHleZjGyrIvbc55t4Q976+Lr2/oklfZf
HKkPC/LCzosvbONptPPXjzcXmgzTg38V079hAhqkdRsnDDLe/v6OTVMnHWk5aSbC7taEVENqIcfZ
P/G+G4VUAnv5m8V+l1Mez4m9SLDAgcNeQuyzGu/tuRtuKlM6eF0eQAs344xgyUVJ1c+1ECwveZL9
Ow+3oG1CLanot1dCO6oRPVWsL4uqQZrwKzqYHDZZXRDZhzZ0xKgQT6NRrAmNrVjOuwbF1wNsIZM2
AcAA82vniKOQE/ToG5uKwsL0/W+XvIqgF2BKhcw0/ufNhGPwK0j3JJhYt2cLACN+1q0xK/htY0mD
+bFnCTvLkk9hBaGTWl4BmC9xXDLJ/r0NhQI16eKuJzx261KMqxwpSNORg/4vJYzH4eylGL1yRcRY
/5OzliRtrBtr75DKYPVMvb9hvRtthtJKa831QJhK2ARdWJhzeSACn3z8tF9MI7J4RxMRWxCG99FT
LTdPh1Il+lV9UUIuSvmG/vOAuBN8RWAObnGDEWDO5V8xnd7fat5DcfRKK+Qs8OhCTZ5tir7ngb5O
IRJIyIeCZAxSy2KJSdqJTT4ccPVz7MZtvW6OcCl2G2keODWU657uU51Ld+XpoWJZlx2/3JY8LhiB
RkSybXpWICMFmc5jHo2JDopmUM8ZET1KFyrZeb3G2xSGLXAmTrYlWsxWLUOSlIetx6m327ml5wUd
dYXgxGaPRGU+8URQ4F7EsOAfXu8QhlnSi+GCQXk1wZH8GrODW6Gnvjx4pEXtom8eLFmRoBtsXxx2
H4Z+pSg2ZQyLNZ4Bne1ahl4y36ZZSZbhJdPdnkoWhQtNqUABm0euFnTQ4FcTfuxwh1swLnn0tRDs
YV1WBRD5BzX1HmrdlTHrDJWajtFpuVuit9ZQVcb05hPGpEFyIeTfh7isiqIbMJEupUzGziJRQaDl
EoByiWu/v07MRXEPwOJWSC1VhnrmDsN5OoWOd+/Gz9QH+5VEksnUw2D20QrtY49+CyGiHzb+GZo1
cKGG28KRgT8iPS7iSmWC1cLOL5HUSRrTJo06CAQ+Wj+o2k2K5tDqT+rDaanPV9sck3NQZLC905vp
D3x58Yq51cj7Q5WFGYfS4Dwll7LBic9ThCphflHEDZtZp+HRK2rAYYTLXY3C0aRhmsZEIYPCqmz0
AxmWEMJcZplQE7cZhqqA3YQQk4fE1j9LYQCrTi/LOKS/SzUnRFwXn3PuHIfEVVTcw0OiAV7YcG0/
SQcRRaR/tiqlrpc/brGdmP294tOFTRrs6QMXeYQCgfwXlOKs3r8THS3TP33hxFf94KyrckYGc8H7
uEQoxGt0jXBfQ4PwNuTmK1W11ynotl/Y8E2T9SS3Pz02EcnPRYWMRDrH2IaAuHpuQ3JoS2Ymlu7a
bH0wfu8G2Io8XZbXs5qn6EyvhmwEqmpaVx5sSOAvJcHuUFBjYV6XmrFxsrAHsqGxSmXyoXVkesR3
gv1YcK4U+vkTP/Ycph73y3MnhVNkmi8YuCyjofLo+ORDCK8QS8OQEKSngjnmemjZ9IM9nnMdXq2M
gINPJT4FFGbMgcf0EK4ZR/gc15mfAyzXb8ZiKe+Y5QGTNxiVV2GM/v9UlnS3yToMzE9bzNgwhQgi
MqhSVY9cYfWV0KfVAAhM4kXVY1+XlZGZB4R4QJZPLXVa4LOab562UZkfxKYHg/KTUKvHl1GMfZBb
P4EpSgD10A4VrPpdT1xUHpxnqXBfmMp2lO/gP984uLi7aNTpGf87XHc9d7HaTYP+sXq62qCL/m6K
V7Kz4IbXO5WPRvyqmEgNGxeSblYgfxA7ePZyuDk541TFmlCsyHp6oLKQ9oQiZDkSffynyreelqVX
8GUbyYv2n1OOVY4NBtuYuULChyREc74jfwwIG4gUCNVXwWRynqmEk5U+SSEi9bslGMd0c2of4Dk4
Sdm1fFvlTBAbdYFjcWbwE9jK7pLc2aO2PQ61uhmjmSSSLsJZCQa8Ji9yeFVzB0A5Nv30GZxI04G1
xkm3iBBLP8OnTS2A3K1WVrESXHrgYQZyHaoYHt4zQF4Ac/F1bFIILGCZg2RCYk9j8XWxCJXhMRNk
aFmNvieopmfEqY6gC82+HnANI+95sHy8UJz48FfKG607try5LBhH+lr/fc7Fq5lfLhdQIRitWPkz
EP2ckqB5yPasFRMJdiDYy2DfuI0K/y3cPr8KDG8HdmOvIJQTanYrDB5ev1h4MEUL73ntXibKm/EX
TOhcFsV6U0g4eEGT3B244iSP8qgcu0mcYp3JSmZhTXFv6fjzlBv9VHoNHK9H8rDCaXbdjk4WH3es
0In4UO6ODxDE489wjLyqTVAgJuY7+sKi4TJMQL2Stf6NwkKXne+cdF0Iok/CYfr/LNKvFO/kJll3
CqLjzsOizPyt1GMqw5GfIYcukmpJsCEc8Pj4Y3ynkw0jZd3S3FgiX8wK71sJATy9o58V5+Bcwvar
8c3rpoWzvJuElTOmEosYpc1r2H/dPFYWASAyiQy+NXr1R/2UYB357JK/fR+ZDrsD+b9rs8Id0174
IYJjfE124Vg8AbXzaUaDv2tYkjPTbZgXz85znX9kTEKKGE2PZcLa991tp5ub+7nr+e1801iBPDIF
2UZrg8ZjWKKHYL4SQZ1rMuVMKQH4FwZRdBinbqZMv8gPIcfJRLppXw/p7B2nkgSHu4W8Euz91GG5
f0WVvB6ve2cGrGGoeIBMiyCw7ShsP/tb4qi+6YPRO5pkfo50x/LWLxaC6lUg0OCSYVHyybjrvsda
n3ZVHfVUwgvJq7l4BNcqCnGro9Wj+bJZHaub1lsIWUTTGFeR96Lc3eUeqj6RYTrPl4flGihehGXP
2S1r/VOtunIkraa2dlTYgRRP1UJA5l7r9KMYNMLebyc00cPX6SgbeNcPnUlUlZqQNQbTFJTPj1/J
n121u+DFZ4qra6S7Err4x9IoQaNE0Lcf0n1Y4JEEZyNlJNLTFI85RMooyNVHKIkwBgrClDZZLs+J
hfgSle7jeMQ4mbUQw5OfD1q4TrXa4lVAXUBwkBjR0H3xl7ywZFwiBPERG6F6SvojU3mi3MGA3KG5
zPRm8fmRBeoZKX9cmnEIX/Phiuf6EXhXOF8nNsb0zqapzyHsTeE9uPlORox4K1wlwu4vut3JBYY/
RDLpYq7japlSs2WecXmmqVrHWLCEWcdz1uCi0xWOUai1Blv9flCOGGM1iMNCuarrtVJoB7i9Biqh
vRFBiEBriFl7YBBBfY25lkQ+4LC+AAJHJg5cAdOXyjVxtfaw7YoIvjlCjNnYMNiqsGyVPvWIy1If
k/63hWWLWltsT2jfmNvZ0v4hJXno6LFNSXhie+lcHUPds85g87Bdg2NSw1rxsZjjmTLlm7kb1E8N
oPO9FQDbABBnaley0lDpqO0T5Q7OzwjiO+HvJMa5RDqCilTdr0+SBSWC2OZ9aga/yieliYmlpTyH
DX5MYhCEvpqFg/o9sy5yBYzhHVHdMpRP+XFq3HwjD5L/cxWQZYy1Yn8zckmIcM8azAoOorLgHAZi
BbeIZUE3u/x+wxWVsm0SsYj6mnBqMAQgc1Qm1vdx7vHqLhVHLcy34f2gVdovi4ox4FOJJsHvR20+
djrUFx9j4t3rVIU45MtySHOBABsvTaR5qIg0fs7dVELhwumwWKNj6E8uKHig7ioeTYFSEY3HAENO
g+I5FxmDXlCQoQWEk+ja3fSrxt4AJpAJN0tAUByzn6RYSbn+OZLMfW6lUT2FYYovzR0rt2ODFu7x
ZyDBg4HBGqtaHyXm5NnWiddNN1xD0xTnq8msbhfkwL5KbsPAQeJDUXRYP1Lt6gbWtTjgGYsArLMP
NlOfExph+bLX6w6H7ZByCdRim7ny+T6scFsm8juqLnBmUtvmOZNFhzeBcLOJmZNmPSSyGKNvHFFz
V4YIocRbyFZPUcCuCQkUw2uvwOkQJC1UvjoKLeALz3YN+Pe3RsP+Q9m5HDuNu1ZXnBXybWF3tYXD
0fgaQulit02PnDNn8nn2g7WYeLqpw4rZ8I0MN/dhwmCkhZkfmf6/OR/k3LoqU9eG3GsonfG0HIbA
9cG3g1XXJnwkFEiU4dWDho7sT9xyN8ZOy4jFK7ylwneB4PHslriCwF0j8NBOQTn8N4eyXUicm5PN
o+AefbZT2gqU6+GUCwi+vki1uIvwLJ/TA68Hdyes9WaxDprYA+hWVuEC1gVkm32XWKe/fZXQt2YT
ELoD1h6duFA1GAHV44YDLZAw959kZpBO2r7rF6itl4FAu9Oh3Q/JHCrEdS3QOe9ygiHbC9n/ZKwr
xncxKR1qZ4auVurTiQBzpddy9jUGVUDTw9mEVgqctHBV7tDmvb3boIMs7HEtvkZ2lnn0Tp+n12/J
E+N6bxZ3xa9sJQ/X8lHWw4mqwwLvgkxjmWSIA2I+wli0pj3uPPoioj8j8HHatxVo+QC1Xa5RWUwo
COFuUpHyUEthNrlp/muYCqjfyD37eRmb3c70oAlwAUzsl4S5qqFKU5pRfQMCf14vaYGE9O9C7mx3
zbJSxEw9LPJfmKugj2Ez3WSxxyagRKTqRDjhq/XUH7DjDD9YPcyoxMlYgDDyFqg9YalaoyKa+bPA
hGCLSz0O5cdzmlXbzM2FRtAV4jx7K9LWNCzmIGQ06EkOT/aQBTPrM1NXnplt6iK6zKUclR2Z76lo
1zKf26SHr/reBYuUGtOey099Ib8PUGudtJbR6kLB0ilNmE0I3Ukx52kkuaQCUrgH51Be4P8L6Ti8
3Mi1Vp4SjonrpMB1WeJOa5oDZmz4LnbXwxsuduA/n5k4Umnv7ZrKiXHSNaJRNB6ZfbsXkKL9rarV
yKziIeSpAMU0eLhJIy4hmyz88GF/jW8XooNUHdYAXnTuJhHuMn8jpjW+UdyJ1lNIe5gg5iD2qZvL
I+zGwIAYujFrb1hx2W84aFjSDGV3BqwCWy8POQKFMWh7INZZ5on+3v4DQuc9Y3BQK7NC5MYYN+Ka
PARdd7VM219Ei8Ch72wUjLZBfgd1Cy+xQrGtog7b9SLRuw13mh2z2GtcusMGLtDp8lQ+zal0v1QH
Xi6BwjSb9vCYGYMvOXt1cRjWowJxR0XDoCf8cg3XhBtOFw4pidVbOaY1Qa6sX9Fy31XYJvv9en8J
uBYwt57Gg8oGLX0z2IkIBwbfKgxUGd2E4RAOUFx4sXecxfYkod+xBspa5k7C+mhKd8MG46Lhf24N
aQd2+4NIKR7imsmZvIlmqG4Bx+hsjh64CAWhp49ScZ1orHadYGdDz0LwPaW/ctcwdS7EtCxnhDuC
loy/Fcs0zi/DRH8zxCOTAyuF2itM3RdQq2Ou9r18DNVOTL/cVYs12vTtblSys6T/iorZVrw/6Vkx
b0+kDoUUpcak7Zq4VM505q07uLz4FH9VD3pgjqXAV2OnwtKVbWZEZA7s9fzQihBufwyJySpb1faM
sKTGZHCj3w4M7Sk8m/5xng8l+IIi2o8dN9AJIiZDHNeR+KfDHxJdW6bcuKbgekb+FKoNoi3rdhE3
v8bAJx7s6zyXMiKGF4zvecHHGwgvXiVg7irnwpOzyAL4y3ghBp7bVFao77Ca9KjAj1CMsgjdgwqq
e/nKZ5wq+ZVWpP8e/oqRlnb2SpTFymp1pxRQDdY4cTzkcT8afuqLL6biecz6dtJ15DHHG2P4jCca
3hp6DjZvp2gzml/5cndVyqSz3fT3QjbEsXO86nW4OtZPhW+VevhGXzk2ou01K80vpya5WUfx0b/x
UgTFNraBFA0NiMHUBQbtM87sVPOYQauRadk+Kt6nUc/fJnAE0YWHK6iWlwXSKV2BoVk974gDmOul
NPM/tU8bQKMS4VKlfYDw/Jbp5bvj0qv67/FNwozV+qTsCESZzSrtVuKEwbhoLy8fk/FsmwB5WrTN
7u3HWBbD7nfJc/sDuzHKUOD+B1GKHBjRP/1wfN+p/NpzE/BQvTXoYGENOB4FF/v1hmwgdO/InrBV
OPrbV7N8VL05EGnBAVL1aPWlvS1zRNHuBSeE7Kw4tILRTMNgzRNmxHWFfe/NsTibjPb2R3bSx87Q
10qbuN6JRk5dLKqajj7SUSaDteXLMjojOX15/oo6A2pViGBQO5b/FXCwoLahaw+WPyyoYuGO6j6j
EWflwvm1Co8AdVgFzOaloQvacmsXqlbWD1USzN6HQn40uAgxXOY/XHQc489j8ZKLEmHPlhIAjGsG
4Xj/mqPMzm0GU3EKLpQKoMqyFz7VB4eKC2jwsnx8Qs5506pqW8/16z/s5Kt7gfj/pv3KidvU1H83
CLL6vyBQVND9B/QPZ/Q9elTjCNr+zytKpjJjwTZrBov/V6Sw4zU23KMMk+e+9c2wA7k8RjQ3StID
trqDg9lj2pbMGysVzvyULtumB2RGtrAFvH7gIBhZg+qK33vlNKYEf8YDmmkIJ3FNMSdKOBoQdPlT
beHQmUycfnlkahXpvpKX6ra0cI/VY5Pu7skfSqekvzEtx6Or462yogGpsEnvYUJ6frpIcPzb3jQ2
SdTPCCL3mK5F7gNEECEqzNeEECSxvj+TJTPLE5rWHxTNPGVMM0zcuV2DYjSXJEDA1C5zimPz5n5R
IxrQPQHiBBnjFHUaOfTGRx5nHixT54EL1GjZ/LQrz8WHcs+AylrjriYfJ3z42iVKGyU7goD/3TtT
PmfnEkpmCGykH2amyOq7pHqPUiOQ7aMep1dasdCg10CWumSfBSJMgL8EFiV7O7l/HwNy/Cdh2WM4
ie2raEiJ5GPYRtSfFmD/TWkInuB50kREBkLWYBgpVtJm2WDKWtEwzGm9GrBpIH6v2rv97iFCP9pl
DeOdnqpoEonQJgfP6tOFYAV8+ksWUckR9k3/zp/mT2tEeR0ap2a8zGJZ+UPCAabuUCf1vQXJTbPo
Tj68Y74nYpETKF4/fxtlpPuBnxWCia9LmcH6C0l9XY39PxDqx1XnWtZfwxcoM20eD3A/1AiGg9qn
mYdCHculCTCC1gm4p8S9ZZP8Yh0s51CzZgdJ6kpx8S2JBlUkCgyLUlepfAqnCraKNRxYFgGAC1LW
8IqRtuJlqpJJsxx19H6Vcm97W2ut/XOiv4KpiuOtND4dqw7k4NcTqzTLJsL0R8Bw3MWM7uYIE/YB
Z8ouTEqewQbQj+RFzg+oBNJq1ULtThwm+wrSFcmZEDV7FNAOU6qBQ5rAyDt2ioKbPLrh3Vfp1bSK
yOPLTBdmv/PzfOp1ZVJWcJMBQpkCv2hIneXwlD8sclC9SKnA+r2ssE+PdFfU1D9ec9whbDh1m70S
WEkzpXXf/UJZ0JwXV4Bri2oGgrkURusAWpKXbFzHlCHvWpAiM7H6jYV5UDr1x7WaJ7APQR/1qDfb
6F5tPEB1L/8BHkyGKnuerBYbSarp5zcvEEG+VzPAukv6CziDEX1LsU1B5V2t5bRzgjS6QD9QUWD6
82/Aae26WiDA7TdlAy6G3Lpf0UQxFLf/SxtntL+kF/UCzHuPaCyFnGGOFi2JWT/I+2fMHFqAQKyB
jOBYdhBZeoUNZGvi9ye266M1Um4DtdsVFBe/QVTdzLEX3ZeJZ1oupMX/bwipsYBw2PltIBtox3gZ
AX3THpT6IWt0V16h/u3OgmSybTCerWrEMO2QtNV7gkboi7x7ju5gEfGMISxdjMabJ0A2MCHYUPtq
6rkqsZSy0Gd+t58nzQGrVCt5OhZeBP21DHIdke4TsegNhzDAhuyENOgJtI9ntPS1zgzVgC2zWdwH
fPvoYMrDWc9eIlV76PMBuRNLnUJNVkLfOlJma+/T1V/+1U+m4rV07Cxz3cbaVVQeCwIfdbfzukYR
oSIHJBZWiFk8Dhx04bnZbs15zbYltNaBLADOBEWYmfY7VD2TOsewkCOyTHyvgsfl5YDlqg7G4Qnw
EKYMvnU80q6AKrrVGaR6DNrXnCxVQNCNRKiPBSm3Cs7GpgO0Ld5dwE2FYJSJccP8ScaR10ZdUfhu
zCACFZXXkmRfW70/HP5/hkuA/iOMgd94r34n0Vml4p1mxj7WzD5ykqm9M7VSbe8r0WHvaQH5n6w6
CAW8B2CR7JEby7xMG/NhqepUrJEf5UAkOmq0/QifjZOiFS9DjxLHxnaywgkUjzf00Oe8PO6yD8ac
1VTr+8G4yfi7BpNf0lU1ukJsm71+144DNcMPCJv5y3ho5h4EVntttuFsnfEJaTw2gWysNihTN3Tq
NoL097a3xPTSkHbESZqhmDVt3WrIzEuVJcJnqfWy28G5+KY8xhd0QPtuWR0lxneD1ufaShTsWyWs
IsxOM8jByFzRKhjmtKYxYiYMclOBJHr3zW+DE40qKehXxMEYjV5E7gRkZVAoSEI8FCCknITPJKlg
Ase4sQAyaS88gtiuBDcTKwy+QWyn9FXwOvEbLnT9hwDZzqu73ib0mknq/t00PBCTnV/oKiBbpSfc
FHN/KyD/q/Razh7Y29XyT6MHeu8RMzEu1QsV7yKKOysa/MFQdEA1ZfUi+opRG31j6tfXXmtYdnhz
ARUuBx//hEMDeEbEUv1OCiXXvXt0YrgalFM4Un7i1a26ZGk9XVicFISXO3TZ3GVAoKFV9B4053pl
Qzk/2itYtwgjyqrHnE187gjD70vzquuIXgfQ499s0K+dqVzIKXSF+NjV//cs+urKB+pcN5462rtL
lb6pZJ4+t9C18VXPOEBq8vacL+koDlbeSqpzWv2RIfZZf+oYqD4J5/waWTtMPWXUAd5DIWB8K01K
f05PsD5+V1f8rBjIo+V9nBuV2wKP0tXfK3+ToTgu2DT82tSpeSaEc5uVSj/yR2O/lrcQ9yn5Cttz
8Pq9aQznm3crK6eOQGZGGMiwNssT6xcGFmpqwg2M9NFgqD28BM3VkUOukG+8eJ1fLxqFOolhOyJC
/dKHdSwe01MwGwwycxih7kaV2MSQFUCjNO+pI3WlT8O5fUTePXG5wwV7Y65W4LP7myB9AsEn/6r/
rdCq7DQ3mz8b5RILZc2E3aDF690DUxerY3yHd9SmoQcmSwBKj1TSUwY3gOvZHsqt84dDNFFneubG
NOCkb4vZzC1SiJZPZrKutKtVuOw6rt7WSzf0L94IuHr+OKoRsqJ0Jq9zDaXGZIyMAcurNUSxBZnh
f2UmJYjah6b+bP3WX5y02ziq3Fmn1hDx1+HaAEZ6evfIaLi+pBJaWyYlS4q4QqcnfLWFSLJuLbCE
c3KbXMMwp97RlJa82AyVo+ZyJL6mbL+JlaWbgjEUkrR3LYrja441RFifAHktUbmOw/zxiUxUC3U5
zdGqRqY1YctKok67bB5ukx33ERIYoSbuw2IibbVcaG+7jLSCiAO6VggJs1uFPfgtONnN7J9qAvW+
gqNhd8ulyiZSHwUkdFAfmhKobuscwdLDek1rlA5rLk/h9O/yMxa4qmQLm5JdVIs3XbHavj3Q+gIq
ifhcn0hN5p9gJs5Gtx86QyPv65pdjgHB2G0h9BZ1P53gKKREKt/ShM638IE4cOkJTM7b/DHQKNDs
yJv1nfwF348MeaMjN1lJhnO898bGJjD/wsZHBZzPtqyGOGAAlj0Pb3mqIabwrwtTBj1oWmkBQ/qM
NQHVzHVoaqbnO3yldqVgcsoCI1Xtc4J5y+iU8kh1Y9FhGyj0aByN5AKcupXmJX3dzOhVSytuXu9u
5FtoPj9j8eTb5orsDREE+1CV6Q5P6DwCWD41F8XMQaxcL443xwzKO2HEFJygGZPi/IjL0/LhTauX
vJS9VPl25jGa/WFqPhGZ+YVssAt2oSEPdLglDLwUOsYPfGXXWCHlociG95MfSa5/9G5n1HyNZvl2
/R4xTC4L+qyOqUI+ZFv3T06EuC4o0gXQJMb5kBvcfgO44+h9CfWZLKcg5FXH7KhfLzXezhqCXQQ5
S06Q2pYRjNpRw+TFbxog06rx6OykxOJ9az9Le4okVDePPAsUhnUCzNtTv45n1UvBo7aHXE7ZamI/
JwkTea6zvqyPEe3KwvsqIpbXOZ73o6y9NYCNja+aFOpxDTdX8tdsxBwgj9EBi+NEdJjXepGomY6/
xaCceCQosecXmhcP7Bgo4yBUhYcRhnvkHhROMeweIm84Gewy/Y1KpRTGPmk0q9Gm3dub9hiHNHvD
tJnp1bKj/NxjCZPXDEuxH5xyuSOIUZLPHczANdAPokqBdwbl0wKfH1tlBums5HSliq4axbh5dVaG
t7FNYixEI7ur8QpvKetY3umnzOOQbiOmx+klH5hBTa3ysBIftgZ+eXsKRLnX7WtGfz0AY1llMgNa
Guq4lcN473fhv6B5zSkRvwqGcswi94thJL4EK4+HUILxweqBcS794iQhr7FqZkN/iTehlGGh4bf+
1TiiJqikNrFZ8S/SKAsleXhb2HSUNBXUmW3BESZiSrTCZcyuSvhHXDImyI+cK58ojfCJ3K5tJ52I
XAGbkc2vbWJNNwAj1U8wAwj2WeowVoRtsH75MTEFFZEKLVlOCgnSei04dHO7Zpt06nlBmXj+BdGA
tQ8wrBNXSOW/hvUHZ52tkIN4RGyjGvLIxV9/wnIDwoswnciyKClhJpY9RNv1ZB3Na6+XJjGEznse
K5qUybLGLkuqHbcH9ZraSumYJlcVykbKrNU61WJezGgjr431uAXnQUQH7TTTgEMl+L0mAc22IYeP
mXH5k/ssDkxAjjKh/xdKxXjoJv02hL0pXRMmtNH+2euytoEQp8ebzaTnd2QeKwNx0pA5uGvqYcw3
PQlZkb/KywngJ8bImhkW89tDvHDIgfgJ4LLgo2QO/7pI9chq3iFygwOJv8OBahTG6AlxZgwO/h/T
hpz3cZORDzYj3MN14UQHJVnBDmiVrhccXKYolzpfMQP7mN2RjaqsgzKUd860GO1lUca2Fdo5tG/6
GuWBv07Un6lw3IuhHqlp282JfrURKxTIQNgxGGlL0VsBEV3VHmLCmXUpMEyloVH59A58E2MdVn2V
+1XFyc0ElBaLO/76oxC+Ze/6gslhoZ7sHNU8nU1eK5wL8NuZLmTwa7HMYooVqUGV98s3eWkLviMz
5poeQuVOzJq7s/g2h9INgkZjWcHQgrSNLSk522RLG9Iz3MaHW+KA+qVuHWjp9MrJDnvM/yUh7wES
7pARqNDgSe2hyKpffZH/uHyEoMaA73SyiUsJs5qV0ghD9A0Vc6loggiY8ZdkcJooHjyDEbSKGGW8
YzZJxP35TWqezoETBiqoEbEwHE6p15wZVjO3WCxPL1oFXz+A7oF6Wl0TxEydKrT8A/gd9o3L7Tfm
vdXLigtSly8SXaib/SuycahmYTgCmS1dt2iTpjoohmb29pXR6fZlWjEXriJCPORHI1dFUIjPgit0
f6wQTe8zS3yTfqr4SUYdlRXyxp0O8Ttb49ux2hqslIpyVQE7n6DA6Xng/esKJirw4l679siMsoV5
Fx0Odflez8yk/MbHuJIGn9C+SGH3KAMARtoRjTdNzySmlGApBHH1ApJKroBlEMFvTP14yH1e6DfV
K7LATT2f9PNGWTJmKQs10tOAbBxgg+/kot9It4gLttBNJIL29QUYQ6TjNZJUt9lEXR4HjyibFMct
arOSv2dizVvQEwb9IFous0Eqh8DXLEysV3cMW5V9LxR4AYb5hBiSpIz6dAz2ldsyJX6w/AOGTNdU
vfhZZA8fB8qL/yehCRewA6tJfRKIKdlAlSVs8WCT4oJa5PFgWCHLu/qtN4qmqAU/lsDJ9mZuKWf/
5MoOAej3kfgDUVy6pie4HBYK1HI2RVLLXsWCBJI7iHEPvP/HOhBf9aUeJSal9tvM+auZ19/hwliO
bXc7F0gDbYQbS+AOKj16GbqdyzT6Yk1Cs6XCxbopaTs8fBTCW688NVy8KquXiiqTO8WNZ0F+MXch
20TgWVcBKyfpRX6/zmoDL3NHWrPYitdyq4hP7DvWPcES17+nUuGWxSdZwU4YD+Q/i1aXejDRPuOa
8r4LJ2MtZAxc+outJAOnUaHR4m4Ne0/XGS85l4uvUzFXQ4Gmiz7nhWQ5QUAEWJJINVLWTqPb9bC2
HL7Dx0S20kVIPj7Zc5RV46KZIZNFxUpS/27nO+uprFIDvVNWNcyAKjhvZ1sk286kuuEchMi5dpuX
3w0PncHFUy0ukG8SvCAv/GLu5V8KMH1wwD1pwpISQq9lQdf15mWVbumKm+RVZRGjOGVIqqeT0mNq
+epkIDW9u29GFoG7MwWdbF2LP4Aaw7SogDr0QeI+HUxqZv/e6MJxD41JHfO0xV3lR5oceC+PRTpM
6jBo5rjZ9ilW/ojzLke4pyCGykFxO6juPYGaob6kwk6Pu8adj6DEAFMAK1DfgmlK2NJd/HekUu8x
P2culQjssJLzUJ2OPh/Dd0GmetIfgAW6wk31lVg189IpsD8nZ8no+6h1R9tygo5qdomwVacXrDZA
cdOKHYbY3qySMuXQ8X1iHCMoejQIBlnwItT9qw6E9o2XBwBP7BO0AZplxJep32M1gZoMG16Ww9GQ
smt7RIihSWRcvzrCjpGh/rZjuzxJ3wac/jhKqdPw1ZODB3d+PL5GAT81th5cqrw0POu7kUlfyhGI
kGw5BccG56W74v/hnsGtRVA1b429qz2/IwzI/ElIuWa/7BqFpWrBLswIt5MBHgilm0fPV8TAqQJ4
+zMz1rtm/gFPPC7tBXgBSDJ2/XvX3VZVsqLw9QwOXw24dmeAMgXht3J+UolIowvqOEsjrMq5qk86
rQrTRNbr37vGbp8novtdhd4Bs+W6PevyFMbVvFYIYzXUEWQslm6wlafjldRlozNc2FIVLLR9douz
fF3Qi+YcogZBGbqyPXFroowDNwtLJ1YsFzib8mBIryToIVnQpgIlJzbfqUJ7MflYWthY7CzFN/P5
Pmjz6icDF/W7MegSG87gRqK41IvcgC1PMfv9x9XItImcm6kX4wJ1aJk5nTUS0JKVLUx0gKG1GqQP
wV4vircjOx7r/OmuU+/dAgt8MBhyRSfx//papudysiOFVig2QXq7ejHFIE0CGVqCrONAesztLEEy
ktrOC4toYpcvI/QnKA7Eglun0TiZivylk+ziOQmlY/vUAOBi+hk0opzLXNG1ENhnrJckXPq8Xivu
pTWVzroj58CSBmj0Xt2HTTAEePrwDDEqarP8t9Dmxa7roeD5XaBXaA+ENNSeXpPI0Nkm6H5AWsWk
IQnreQ2aUj5mTFLk0RID3tf/KOibg1w0c5RZsOW3lKdi/oxqB+JI/tvE5ZOGB3sqR2k1UUhfvNhL
VNdVjuQSj8p14Inz5EI8EWJgodnVEZA/nszCVXnUTo09NVf/Q5Rmmzl+6kqxf0LJOi607GW4vzr4
Mu+1fVRzcQc2q3m6ubPgIxVN1LIOv6ogiuyfexsTkQ4xH4v9pnDeASV8DqV1/UocRBpUNKQJtyfh
q7f/cwWhDB7vnK0a8jU/+EZPUct7MkXvxwHwgOUYjo96AZUUnT7q7Qy7pMAZ0GjvK8p8GALsYLfy
w3dibhEveuSiyM4HpfBday9WUMNLBudRMa1hj6k1+eDZQEHczBj7cW2k+KH2N2lS3dPabhjAWdrN
YO30gXUlXqqAZbLKWqrsnnRfuu6fwak1QwdG7naaq5GLbtZvR4XDi07xnV7JZnuQ3z/kwVOdkSKb
Q4qy69ArYN+cYZFsYG93XAMiS+Sxj9NsyyuFQUX8RybHD5bYcknpEMZFU9YRCIqJ9AYY9iDQWQ1M
/Q/Ll4pjHo4SE/reTfjEwkvbcB/+Qv5EJoAJaqwDlmK0wf8P7YjimpPNByPWnNJ59XmqRGjIFZcp
L5g2Yy5c/gv+yWQvctXlfPm6sRgPnKcxYzWVZ5+6p66RPTgWcZeiaqcP6ufbivyrwL1lN89008NJ
wWKrPDjLF3DDLUqh3Im44VD7JZwVIL9Gh5XuVCkIjMYyX0f2C1JduypcHy9dhkz+czkuLVZBiMjB
oeZ6XqFW7oEfAJ06Stm7SdL9vEIJdLc4DUfCIbE4YZfVbMN2j2nwi0MFUmYU5ciCAZBdwTXDPPgm
90krAOUFJICbEAqLbD7snfxGbudRVjMFK1uOzeF8xw2rLkfwMMtrnRGBKSoFCAW3ffamXGBd6Z3G
gB+pGge2eftFaIMgH0+cKaW8wQp2QYzjNm71FOIrCsRttxEMhuKPIVcTIb4ro7QzSlumvuJJ5/1B
vN+jTb3zmE5ufQstEKKkMJessaCS1yLaL/ei9Es5RbZlkDF9J4MHeVz38J6Bs6zBngh9veo5LfYA
XB6/aIL3AsVczc5CQ6cO5qsbuEhYugKH7VB668qdWwu63d+724TqIhJnYJUdapKXFHO4zY9C7rO8
/oTSJImS6JqwPP6kogMZTJvuP8NfmsbC8aApWy4zddOE54vxYy1DFWJzcbdTRygM/n9Fc15sHMLl
JfPvCOGYMS6/thG+SdeL9xvjSMt0QlfiAsXABOKvk65MT9hzflOboEd4cisFioq4UNn9yCH6N9Tn
vl15YD+ms+Q7fgKXVGofNxxG5ym+28qvpr/VSvqaHKyeCppNe8gyi/vfwLjwzAi5XXXPaS+SrP++
uOFYejV3wCmSHo2QyemtlrW80tLbnNcOaJwen9L+H8/bQfJE3OqjyaQwLSb/qxMs1/1eyVA8nWDh
PsRt9sK92Rs8+NcYrI+kTdKMCRXq3BlR7/CDjrUssXNOFxjEqO8KACmCMg6BydGW+TA9qqFmX38x
fuK/qQPNH8+wozP4CzerMmzNONPIeOGZLuzOossvOSsNK2KUqjNIGbcfv0c2tO4m7bBUKO5D3dss
Ho1hR0n2A7jUzYfmEYO3T8/YuorNEbqK/4j/rDimPaOKd7DXv4F37znD0IJOyjGKwCaxE9OP80iX
Nt2yjjsYJfhZFoQJI+eNEMF5fwtnhmQI9w6B0FfWNJRT0PuQ/28am+sG7MJiNwTR+yDTLmHXYmNM
iqRs0N9AGJhHQUT4p8N1IMJG/mkKZLvhjS59jtj4MQAa0ZEquBbisFK3yUa/hSHAfTYfucxTRXpT
e7JJBS1sI5f4xaMnZ0jssxlK6Ud5WMuZT6J0DiaA5r5v9wa0HkvcI467sZnWoHulv7wr+pIbqkXL
bMxidHu/kHISpvj5Y+cKfDfRKKbwq3y4WFoTMKYVFlyWULOikbLEujrCjDVXgJNRsB2oo/d0aPAS
kHgqZrMq0/QIuF/kiaKNACUGQltvFoUUEj6npLpWXDR1kJlvXoX3WIZiTDFOuo/aUxBmAFyBfRbL
xDov5spRn1Q5JkJOYdJcb91GyKeLASXyRz2Otz1ZZ777ucA9+B0d4i+Gi4YjRd4IUCSFHPSSH9R1
ZUFFmrW/fd5MqRakk5gj0mcXrrHlt/r2fAe8nMvnYwZ/DGrMVrzGlXmzOaRhWCRILHLf+rUlcyXK
C+dsDYLLyjbLkE5g1kraTsVRdHiwExGh04zAPZwO8jLRlzvaNwZlx8v9sujF+oK2QBFddaj72RKH
Gs5TL0AwvMXSqp6WmQpVKQ914o/5SLNQ06fTebatbDA9RYBAhFSM1qS6WOcblKRKmfjgcr7N/HgC
XrRP+f65EWa6/IJn9H9OWmNvneBm78PZO+bulC187gz0S8xyidGyAE0xNv1xg2kH7fDx9HgknSIr
oSuLtJNBWXtT/o3mFp9F4TXMohMVpUY6BTAicq95600/EbvVEml7Hfq0sMecuyK5lN5y8Vm1EALy
I9aZBgJlajgSHQMOWjhcrSEuyyE5/v4YyHswMeM21xX7MgytFFbLwmDjmBpsYAFaF7UbCYz4NqYI
G6IBSurpgLeEiTAK8NnhCfiD2zwiL4qbhELQeEB7L/GKSMozRgtDtRhgGmmeQjngiNR8SYN/UpQs
Fek1IqcJVXnZ3/BRYKVQNp6mgLq416nZBUWJqkE/Q6l6E4K+wxLgXpXjWyfTdQwb9C+8g83BpCzc
ZRTATPyrKtRu3sE7MVedO3Dvz+e3jTCyYbyFxGATjSNtP2LmLcBQVaOXxexVl2R/Wc/A75H4XGqO
CEZ2D3RiMVkeGNdcnWOdIUUWHBlWumrr6Axpgon575q3ub3Kui016lMnTEOesRhNL6javvd1M0E8
pSsxa/dk5C2PG1J2m1aNqrhdvgcTdPuZy0Oh/0ziu7TO3vgM3JMJF2q8DZlQymJkjXrII4MmVeRQ
QQW0oBEgLf+yJDMeuIqdUZe2igUEv8/DlgSYKKQSktxky9be/4WMH1smijqKMe1JhXf6gKlDeoOP
SuG01axYhRCDK49b8RzVtxd2E2NdZi3w00oRUZeYPsW5ZYT8nTph6fA3uz9px2hp7FE9sfWOdYr5
pCMKOU7WVFcUjZfPl7LFxrxJk0qhGa3nE62uPs3KRrbuRRYnhkcp506PyyYkefxY5NqWofPHTxi0
kpPM80Q2kHz6unXfa2S9Vuah3jhRTFMMN9u2XJVeRaJWNCtj2Ro1WU1WHp0fAhGYjx26X1KJ739U
zu3UBxkF6GQ0/axrw95XhlSVbYs1PCviQ74UY3y9uk2hZxbfEFNGZP2OnisUvXHP5DTfQjWov/Rg
p40kCf2av3U8jMq3Z/iH15jJA66LQLCfIUVuwf1yeQp+2O+OTCT1odZNPnDhOjERdONfyUZsJ/4K
DgIHogfHRMP2FBqoUPKaTwZelNLqV/d0QN8H6R2PU7Y+fpTb6EgPsyHTmhUC8rqW9b+sLLWb3zzB
NXWazeIeMdZT3Eomg2Xxlgt0YOajYYMerQkHA8bx1GpHY2H/BrNhi7ouzTuVRaIn2mUDJ1K7gC2u
zZAzjCQZkBY+e4uz461iT3eibU6GPPJkvUeB0YIs7etTNI0nhDHI5kvdJNVBgaLHsnj5C6x0PuG5
Ry7+8YmDS4EeH+cg7fT8GbtE50kZhh12mTXxfrSnpiQrmAQl03HtsFtryGGnl6w2ygFW9DPoIBzz
Js2ujYE4iPtpBwOv+W44C40iSqZzbtE+Sb6lGkI4YRG99r9fm9D/wJH4zvwIkkPgMC0k5Mc3hTso
hfSS+sep8s8BWYj0BcavftE79tiIMSrJ8icYYXJ++NOwnHxqOMa4V01/QRU3h4Cd4nL9YcMkWGZs
woUhxPI50avfHdnL2lJcTd4D25wtCUGe7hvyvg3BTkTRK6cYCnfoItNYpUkMfvFm++bY1+rFyA0+
uBBYpX4068KV2uPH0aF751KOtpE9jMEKnyEtpGYBeLw2xaQJEl45R1pnlzaVZEhuswQWsQrCrgXp
1x54k51Ab7MRtisu2ilS5ZqFWsc3DeWnCIY/9W3XMVwjDNj58JX9F0DGf93VT4rq//G20/TCszIq
uhdsjCnwybQYeQ1CF0mfYCS3UimM8JE+y2Ic5z+hBOi0/9W5pYEUdhGJVnmfnN1GrFMQoLbJIQix
jXy2O1lLxqokwLF+50vq3+oASO3iAoa6RzfZx60ljy7bv7W/XUeNJEclyRqpo+En9FcACjH+vzyG
fWZyel+vZQlbyI3SCihA590wlls6Zf2o0vkrqzbT9tB7n86BRBXwj3ncG/0JI+AwRxZb3H3vmybQ
9VeKksTRm/3n+Uye9h6rfy3su9ZLskEii0X8tjzpu7RSc//ROIQZ7bE1YqIy7kacszG/n5iW9OLR
e2LEiD6G1YllZ2jn6MNRag6oGnNJsz0H1F0yJs1ULJSfhXzCuEc6znGXKyNp3ddsMJYfiBarWgNh
vQEb+8DBN0SImSK6Rm76V8Fd289G3lUibE0h1tRYFu0w9rdpu8JstK0HLxxt7u4keTLmK57Smk9G
a6URH96FY+vZEc3bJTB6CGw3GWAc5lPwtcNyxoizcgecFe++AulkHvItw6rzqZ8w/6Tb/5c89TCo
RjAhMMO69PkH4BwctlGO1FTIFlIi/l3IfQRQLRcDVr1mbJjtYUbjJAs4vXERMP3JyOMqGqlfHMzy
L7mruxTN2UweBLTMkrfzf5Fw85GhMLy40JlnxGxJqg6nYls/fVAKcifj0S+kDXnYxEicWJ2kKIvK
a/UyffsxpDPUHSQmYorQVCdcMjKGwxBOd6KUSIqgYY1zRdavnilA1ZyuuhnGvdZbZJpYqnmjJkGa
l4TnQuqS4c7jsLDyqahhCZ7DGeygFDTTedYQZ6Z9lcqeUwIdwRV//XFMEpM0FN5LP5sLCfYM02ic
+v7Jwo9exs2wQppCgJyE7wOckjIM+5DTLPIIQOQylLB7oLwGa0sQ96EuZlXpBar/jqekm+iD5QAA
tdciqYzKPqIJx3BtvxrA03LmffozkecbwLNoq4dTKfE13z0gMnwOkGHJdNJKJkRGeE/bXq3uRYZQ
owwPv5kzXm4sPwQI5xSIYlIzE6qkL9HN0EOBi49mp+KW4GKze6K52rayVzmBFqfhAylQQjSDMNyx
9xL59qmpwpd3pplHfMAJZ7qEdcSKVV4ExMg8Bp1F0YuKaLZX4WL5/CNtLqI8FSVbDWBIWZi8GXRO
g2VCHWBYTyhIJHWpqKXvlhmFp+gLjTR38S/DoqTQYOwDqUD3Mk8yJE02DGSRTdqnMXKWZCS1ijQF
JIXNk2qmvqT9YMsLG222hWNud1w6rv+lW6UekAsr1Pt+jmfufFGhigSNZ4LiQVNZJfROlnzOh/tq
MAFxVKEzOyGUxvEuovmzsMSb4yIqYIOEVlYmzldwWxc/NThKAHjD2gO0iaOetq0meskG0EjcIlyc
Je1Ywgf89DLcU+pI94DupmOhJblU2a8LLFIOJgLZ906bH7OE0EX3YbawT3HRvNKvTVgvOgoMmqr9
aYPZp1D4DU9NzcoOnLyeMfYokEw5RPKAK+Gy/PNNphBASUrEPOyOT+pt8virP/VduiK55u9YZHHw
x+doMwPT2zZy1OfwdvWl+zi5BHiUIVTZXstSAFVLBQ2scKBppskYlpUwj56ZXdbvCFIhxacbwyxL
YNr/3dcrbTEqNUKmu8kcbB26gyA6V1rCanKH2ECLyCc4QFAufM762vxgo6PyDFQhH7frSQJJshcj
LnwvHgHKMkyqBtxd11xaQcslGQvkV6Fn8fbv7tn2MNsyX2EzT4SjAdCpYMnEyakLvjd1sQfOxL5D
S5uaap0D7pM1Mszvl7KIG2UVIKcdM8BHzcASmK/gzxikGn6+Aulm303/MtSY0rDKoSf3q/DR56VS
c96vslknrTkFCF6YcJwclP4x63Vhskvzhyz8311t5RX1Ptb+LsfpAM/S5uNcOl+Zgy29kpWcEVjJ
yUYlUSg8XqW0835stpsVKufMLcUyJ+7DwiWIw06G4lWWwhNQtGeahGvSVd37dqe9fzmxJJKlfQ5J
PMv2IwMK2XZ6BIQUZl0Ma0CflO5fzl+0Rq3bBeTlUl1GalEDFHOW0M1seTeW59/sG6MhoQmTQ1xZ
5KFLpfbDwTsDCJ5TKCJJC2W19iAgOcMS2yOBOPiFsI2ETPfUrQEXdSF9GEnVCkbXWXxXZRrgOfGx
tgByE1qxKYH0C5Kby5HWIJrGZzENxkD0jbHtFS+4LZU8Y4KFYmGkrmCWJv9kGI020HVEaAJ+lHKJ
OyJ9b+aKFctQVzIBeNnEZhKcpkPSW0RLwlMQR+CFbfVIOUFdQ5Qmzp6puKV2clIle0DN2pYp3maY
lOAH7U5c/DiwHCPx9ZghnmNBYTh1eV1JGQesJ4ijryvbuhhzM1NIUsCOs/wWeUvx88tQ2d1VsRum
F5wHr7V8D1kxv6XwdoAQ99NjTzYViHdbmCM7SjOVXl9/+h2jW5wMn0U2aQ4Ln5wuWOstQI2QyW6N
Uvt6bFyQU3XaCE/Ka4F4w9IZ3RtgiAzDxdr6evr+Kb3z/kZ1qsrDRLAyL5FsDC8Lgk8ZuqchG5hB
9o59k6GB0O64UbyImRTaIXEm9hutCg7cUMmY/IkYLSHBqyBLTgdRuJzrYwRJGq+J+gWtTmfoPRVh
m0hkpYJgEsKufOUJpnRqtw/L5aSnkJFNe8nWLKWrwjw4OiBkzkfX91fLBJPMQ879nQbMR4OVpaIu
LzCbtBzdSrkTRgXdrbRHb6WKEXOabvfUOw3YemQ2TRbRtbyrGgLtTGlJr3RBX0EBtNic1G27P+Om
sACVAXoXyVPRH6YYZa0nXooso2c9aOj2eKXdxgkQ/FeoUcplwzsfKsSvN+OBoJ/YwQn67U+ii+UG
JS54WLaA1GpUxIav/LCyNbSK0goSuQ2FISl4EG+VhIKKU8XED/eQirub7takXMPJeT/5dvk2eMWt
HEJxI1RYilSbRbcXrm2cATz/N9U26Usu2pWD/1gDQYK5xNEpH6I2n8qCxuP+DOZXT8YPDEEgxYIe
eFsSEInkFo+sza0CAp3JdDdEjBpM7w6hcylx/1qNPQnydXPe8dsBYied3gyWtbdRr70ALYk1mljA
git8odrYE5lzJzKipN22aSTEwcGmLPXv+oM2HmefJ/vVvJrQ3c0d5ApJhIe10M7W1hgZEjvfERz2
xBVpoE/etK4WOPPxii7Jo8CRWkQjbCnrlV6qrgWOLQQOSCQ9ZGLNC0N6CoKgasFrDWJB7h4bec+A
YZ8OWCjz/91O1a6IV/th0Br4P0yjO4Vs+cB77eTIdG+PWNgPRt1UMIWjOEXcWvKslMvOT8tsdFZt
UeIy/dydzG9to8pq+RW8budKNXa+mMkztlriTqh1aNZCA20ELL/oxvk6evMjXCTNP1Agq+Fbxzx1
IGAHdGoHnawhublr/syelT4Xtf2ZaU1Y2Y4UtVjRPqZNumB8XBg2RMDQNUf3m8ZaWoNtkZUfveiz
aV4H5RLVIdUQbXrPjK+J3u6avLOKnFFOdQrVDcqrGu7UOXBMyGDdeezON7sCSBituIeWf/rBXnlU
NM572NnbQR9MVAB2o0z6ow/oAJpOFB0iUbGA9PnVuf/5ITWWcrlfM3ec6gK1Ti430SLFwuouWdwa
Lfrgm8KdUkLsHvtXosYHtYuGbwxqUuNSmfmBp0ZyKHwM9jNYyJAfeHmVeR64e2Gk/0QoLgLFBoJS
bICJCqxzxlYk+Yk3x5uHJYCg7bmysRhOuGRawsBL3Hf4vZHQ5PGRy9M0zhxhlXQtblIGQztlajJ6
+fNCzK6a+MvrcYZFOp7iPgudKobTEqUzLR9LmW0Orhha0mIXQ+xYvCmaA1D9vB2yGEiyUj+us047
yBjj0wZ3Cw8XbRcAjf4YHTxNEnFcK0V7DxpZmT44vdJMQPtf6+u23W0jZVaYkz7RMvtwQBGSarmR
mIo20Cf0Prej+AkbJsen3JTPNY4tGyIzeva75Y1XMdJRfdgMRgyekaB2qNGEtouG0o2ICIxcR778
S3dm0dG10Kw/l1E9ycUN0v+mmpaJSbMezmbqZt9wpbJP4fB2FJIOIIHsLgfwGPdf0idpthg/7HXx
pJXmv0poXAUN/pHU9azUmZq9ihljo7pTmkfdHQxzRksi+QJQ1E5bD4L+aHDJq6LMAN+ZRuc1VGEY
6e/B9/tsKsTlNgoIjLv2QmcsoCqXm6QyUeVhaJMKC5Xa7MZPvAzjjJZMGAkz7S2XF+1NCl7YrRHm
C4AUGoFzjBmPGuT/DgkLZNkMyRQKBpzuxod5VFW1FaOss/JwdNf2R+iqT01OATXQdwA3q04oiEX0
t2GbkQ799Tqr3mumCmnYOcSA6aH4MpI1UNCRzejpvLe1OvhRDglpmdf8KVc7OPxjpWj9Xs21RIqF
VMah8isbr/nDu3Se11c/VyaH9jfLGaRqI0KBkG1g9bNi4OV1zw/SgNeVdJ6GEQz4bdNdICz6jhd5
bJj/IokCBYK5N0FbpQYehP+Ui3kAN5bSMKkqTXYEhDXhcPp5XK85O87uTohpshU/nV9edc9UYLCu
XMvNr6idvVVqJSJaQYPvKKfzc5G3KL435Y716T++bHbvbIFinXs2+s/JEXxUeBp5F8QvDcV5xQHM
WeEcLypor3B3trvryyzqmlA+HE9dfL3KZYgBzKa+Jv58ELSmqfrkv0OcLLy86Y8RiqC/A4RS/S+i
ALjESHsvphwdsuYUGlgkVkhEQRKtUv9Agvb3i7A55Q1GqwK0ts1BHApnvO9FUvupTJFvct3/4m/t
m6oPF54S/BhvMETESPHlO5HPKLo79EUFvRTUa2Zys9a4orT/+E4dIX+/PZyUL6h6gxanv5ehHE1O
oWSimCd0GB8KpyG3f2FW5E4v/29qahS405AOIp7+tILdWoO6PQhRF7FJBdscArbsN2axlqwBxYEI
1d4MVYCFfe4ZBlSF+TTHwxw1HhZMRCCxNYzDUriK3n7ezUUCOWUR/lpbfCsLR6+Ad7r8o1ZPJOK0
p7pKI+2dts6X7d4ZGdakWc8FEAngWpwB8btYJkob+S47uYbc9Qa8YU0MJcneqmHy30o9AXhBMx6i
A83xMdJam45s6IrfYpgH2/PjQs364XOVnmmN0+y5DsuREXnEuX0DaY7K/zFUKhtbiCbVlT/Xq8n0
JryVhmJ9KD+K3oF3E9cYoJ60/C8WtEsfEW+TH24Uhx0NCkKe2jRUGlik9sP1w3LFG/u8OpFPV/u2
xL6WPJ+TffBcsr31nQibiV1+YqPqopYBV2dO4OIOJB+J7gbTlxPORlmC2KzFvf1nBWfves4XRHqW
UcQ7Xm3ThjQZltWkTFjPCVf/vhStkUuFrWCtUkaQuX9a/aLh67tUZYN+PR/rPRWWtb+nMqJLmORu
uaQHpSPTEHz5jWGr0O0TO/2svMLGa4k0vVp1jtZJq+Ua7KE2Qv7HmDNkVrERY7aKjs5RFRi8OUjs
HEbtoBKeNEuWNF765ozAkH9l38aVizLZOC+en+WtiqrAulnxUneY/Dz5wcPzDGFvcsxKK/8N5NmX
vKoEVhryc+bPiS5DrIEmMk7L2v//tdsgwG7dPbhCXDXXywxzblBguSI8nYauaCFPDS58myz9EHxe
GIAwYBz5WBTYpO4gufFkWVTbfAQ3q3m8aMtbtlHS4fs4lkxd53J0GMBNluAlS3Z9nQUvU61/7wPn
MZJhrs5zwgajd8oYH3z0/J+f4hvuKTgzokmbJQtGE5mZ2DHD/qp4PPGoMRssJCcHG66F1PkVl7EK
zZO6DBjAgqRyL6UClbRT4c18vB8NkqN+KhTgg5fy5qZZAUsl3AbeAGflMxTP9bCXs9MGNibiMaSs
4B2TwREYOz6I4xVActNVGlkR0f6ehxWfhbJqYrZ72LND4ljBc970n7t73ynRnY+nICJKSwQqtiPG
oXLfijk+iT80pAJZ1kJ46xS56Xi9mGxk1kXmHbaQzeU8TXJpO0x/qSKfuaancEoxOYzpWPAACm1G
MXkZRDVywdWaO/P8FiyyrQ3ouGoXg5Im+gbpBFKnwpEz6WcCQqTI+tAVl+PhP3ynoCTolPCFE2LF
2iWoksW4vICD4K3yH3uXjgaOzDZY2YHuAEiMStqdzNPOQQ716PuuZTS/OjiIBkiXwfwSTLzTPtJU
c3CbCoTJ8Tbrl43FAXIqIqS3LTDgRNEyNrCVIYLr1ACRrMQglWEVNEXjhIU1ChoKfeAFDz3nxHNc
xITH+IikwJWwbWSezhDczlAYYL3x/iKnVPLJgwBz+4fkXNkDO7+ymZjDSX5FDY9GJ5nMf2OHLr5o
JXM6W0yEFRBQtGPfmTHLhPsAGqztUhJhILdtL37lcHWhOIEFFnhXkACQ4a0FtTC7rPZFaxzLOued
96u9X361drPbiO+urk+AypAqUgVlHr0ByBvsPeKdBWheA/MovXA2pCNNgK9PAA6uJTQXUEn79C8i
Hsca6i/aQfNi0xrcNHXVHigypp4FrxqS8hHW5bAIhJMWsevRsmLOxCYbrvjN9V+9zipoWvDqqHsh
/vpvEr65jqV0KynFvFl6+75wkbrnyBM+VOm5UAmw5acISohiPVKAd3DZWfibq8uGtHpYO/kIuUGU
nErkgPwY1G9Kh1U+0WiBmXId1CyvKvNMCByBCoZAFVuGH8Nt0dX18OGiOUiOl6A33Y2anJ6bdX3e
DfRG2jlWSL4eSLKYRds+rNCKyP36L4PK/MhtPDH+8ONgCk+oO1ncKze8Q+4I++oc3TbmxlaZON5y
lLlkc6dArXF8bMtG4C3svEO95fn5/o9dxQ9kpR2T0fGYZfExF3aAqf2fanNgOfnb0zENMTponfyL
hh4i73OjuuZj4/LKnrQ+OWqVn4Eg4uSy/MNeiAmXZ7M3XGvuJrV76m/PWer8gGYkpEE8KnxlnNEn
dOCU4ITXfiIJ2PXYNSaVWcntx3u/y33Zj/0Hfdt3FWqeKXzQu3u0RY4UXjkYUBfztYaLSTJBQbq3
rmOMpOJK7Q/768bGi2G+EvOJcKvUIqaIZuYRlNNGLkyWOitBY4DylBIBB3YNRDPMDZU1eCdTva+r
OtShlwbTR92Mij3WmK0YndRjM9RHOea+SPC44F1Jf2cGiNogpNKjZKLr3GuMfows3+cLE76BCiQ+
bbXMgzyyAScKA7Dv5uuVB1A8xRNYCWcIwEM3ftvu9z9PJLEywBWGfQe9sjc/1a4Axi1IZJGbLRTU
lu4nCF/MPjnjJGDsB7tqzUqQ4GmCN75dP985ryVJ5jPs/poBzLYotoN/5BaQe4qpVqkG6/EfiEH3
o3jh3YKj2o3izXcBKH476QjgcbLhStzFr31rvCEHGcNQEkVTvHRa7I5LJqlrfL6yQ/7P0vOX6sgc
hjcvDhc/FoP5GjTXT/glVDuXF8joNb6X7riSB1/L/QhltsXdzXu/mAx7/aSHlZIw/rZ2mBTj8M8n
L6++eolfsSeyYXa8LyWb0ewhYNXS3hFL/axQH4ZqGa6MSZLtZzMhxgFKa5FwcP2+aJp0x5pMM0FV
fDDG44Aajak8YKjMGa1d+rKNmr6p/+C9JyaUHzjBr7NK8Ozv3hGTfZ3fJv03EUnRjLMLPygk24Gb
Dj8He2DQbdyFS8qh7Iw8caBk0FanfJs2bMXVQYQ+THqHSQzwFYZxDBcn6MEC88bgYQKHfrsvPrHk
G5XILm0yNGl18Dvnh5fKMJDkpP/R5cYQXfmIDYKjian03I7h3Bw5zwIh6TarKAGl6VXncKkMNqBI
fb17GjKhqp/KsDQW6aCHls+P/kOK/sEhTS5wwfvyFdKuUuE9RnLHDVYymCYYhYDFhmWJtm5zqTNi
ha+RV3/zqRBho03WAbDD6p6GiYQ6D7EzD8UJisigVtX0KpgB/gxA/P/Y893UJcBQm/zZ0frB/VYZ
xua9wHHL3NKueYqT1fwCiySSv4+EzH5o6aLstM1rrVsNkHNDacmaEdBEOZhmTPdvhjMBIE73H9vA
EvCuTaY++FtY6mvZvLqTAw3e1OiVuVJzrSsJbJ+GZqKgGYPwTRx/mum5zEwBu0jqTu/xn1sjJQ8D
Y08Y6uTIfcIVFFqy2g2ENTAvaXPuoW81uKRT4YTpEQtB5Oj/tWD3FIHnY7aKCwKONvyJeV6W6OaS
mFbviqnfRYrVs0T71y9bZWwBcwbpzrQuk7nL+NOJHu5ZBti/On84GEj6QLSx2LPiF1O8JUOP3hCN
HY3hNGXVJJQ1bRLh/08Q2tBp+kpupaEb7YSNATTpaHEvKewZoTlDGw19XhYAcLIzXv5IBVCAdYqG
F8w+5KQLKS0KTd5V5fKxe698AuS2a1MXMnaSQ3FI3g2eNlwKPY91K0EFlHiCowTW5Yx7mF/xQmjL
qOZJ1piPHAKb7/SGr1yBr2sVutee0msDaadZIn0vY57PDKOZIQxNZpazkIQeAJzrH0CD+lj3S1gA
kydEUDsRr0SARiJu39YuLWHVZJtZqxd6kZMDVRQ+Dl+ewAsG9IrWder52YURTW2pKFNnv/p7VjZz
Ps1VjAPZKrA0efhX1vbCF4eb31BhOuY7U39kyK5V6OkKetEJOZz7iJpb0TWCUkTKtypPKgfVsx7p
/lh1BV8smoHoYd7p6csINNwEwGQdmHVFS+R3CRAmbYsvAFq/vi4hBLOFQherhh6+08EwfgSfXDhS
D07mrCdjRqYXuneyie88wFv0kvcpufdo1uHK44FNZr51mSk8PIo8+mRzqUMdh72ZkAOiRZBqZeoO
cg0o/uXdJkf4nqTFS1HRqXE596e6gvaBf1ebt3QxQ3QO4SThYji60fnKw2zSH+Etm4YNcI82g8i3
2yJRCl93YZmvrn3NyUZQaSnVid+pNHGRTso6vgFyR6W2/vgoWcKdOOvyIEXgC6cpg68qMHW9Veo+
pwFppXRIUaZiUy5/hXgoGD+hPyee4LDDZYsW6qczdPLwUArZxwAn9/ZhwKUhOGkf4/vFSwEwB6Ku
A5/H3dAHBp33iBfsgKdq5i0ElSikqoeXSxJAFrFo2Ca8T8GxfKGrfHeE13mJJTZHWO4vFoNMz0v1
LKy0Cm812UutR4kSiz11yc3atv9QNjUiYdkUktbwps4V/QGp7hFOELEVT0aTkth+JeypGKhoHol0
Tkcq8fMRz/aOAiLa9UnBNEFWXVB98lBCJFc69iF04P1QYv/itEj9BKu8lfbaJhqr01Lw/W/IFzQT
VasNYSPRZPErYAsQroIuJmF1PPtdkm/pgeNklndcuvhZBZ5NfU1NGN0isECK/oC4USa0YBH8o4Z4
w7CACSw1tHeesQgejAUZn9bT5LB53nBwHCZMCaXUQJDjMYKJ3e+2J99EqX8yqI8M5OFgj9dNUYDM
Y+GDoPcoW2SItR2p9RxVvB1jRpO7oIohJvV0BJeR5wjvI/pxul2RpdnMquSJ29Hke7UbM1ucZDMo
/fGN4JmsldenXTSwXFinJ5k5xSAahk0cCDbf/qHlisA6XVgl2lMYN8+yTGvkqQmiiLhUOKBtbzhN
jRKpAp9naS66b/ZrxbKJteT7pg+H7MRJJ1wCOtKjfqu+0Kc58BqUCULZXZZASXbvTnnRfC5KoU+U
SgPeThX9t2sLG/SiI3ksXH9PHoXnru2HelGLUBvY63aHGYmiEfXl8eYGl3jdwhA877L9NOuasjA3
hYTXYaf6B7PYmM7FmvF9FfqligRNP6EedM076vu7mTzXFTxAVMGaA+NEkQ4A5MPtAh6gsBEq1MiI
8Y8JBP3++yJpdLG2WQ1kqqJK86sOG7KySuhJvQxS6GWvfMq7Wn8dbXbnFVUMYw66xN1N+j0B8s/t
Yd7WTYst6jJoKZSnfMVbHPHJ3Oyb6ITXaDTC87s6tXIHicB/R969HlEu6Bwp1b+2lFpdzKgdoEob
sQvZxiEUZLZaVFttig2jLS1Gz3t5YBZpKGPl1QYeUJFrjXDT0EzS96KOj1ErhsOesEmr0g8ocqQK
hQ9riJggPMXz6FlPECcad1CeQ03QzRbdNsQo0hgy1yBYnelOMuxI3PUEfHHf5Wh8cARsOV7lKkyL
xi8m0kVvVXEEaLW8Tp8jELBrm2vtrMNF8u1BXFqtl3jdwQIcJba85dAbo/kVqKCBbK+0zH+FbyS6
RD1HiV8FdKEN999LQSciNcyzHYBnImPgHn/0+a72i/2KRNzTZqvpe6BN4Zm+DeIWuCh3TzVreZIj
SuU1lL/DRy6u9f6FUAay23tBTXQ8MzYG3p/ncl8dmfXb5FMHFLsd0AYxtqpjjSOaOXzddh41JVNc
1Ru8Yn+P5gB16RSyshoj4HM6QjZoNOR5jpU8TDXeUb0S3V4kQjrKHtCtQojF0KYxbhHn64UkklgD
/uSAo7XIbfuTdqgoSEPymdWOwInRUn/8ANG1NUaxdNsKprfm+nbfb68bYKpowYCNNbHcikdy9iZm
DQVUVnjyFQG1hXmwlwrglofyJobeeB1J95rxipvvJAERanbfb7VbO+nKENHF3R5H2nbQnaEyXzNG
IHfDVqrAkmS2rvkvUrkGJlugEICTx/SE7POvuXIefuUoBxYmQbLB4W0Gikc4ovH63W0aR1tlrz/5
kPsWZytYOeJx+dYZyZHXAD3cvUEF8XtQbFt1oOxNpRVoQRghIp+szPqboLdPzFrWgCmpUOpe3aDn
oUkqwfWNjtBbJAtnkcKvhtm6CiLIjIGiIIpeARm9IScVph8mM7AhZTlFL53dUS4rA6Q7DK26dS5T
ZcwFSgDtNnfIPah2EHwZmn1K9mW6+F4b9wkWIdmrXCBJgeZFUcLYqMnFEQ10kB+obJ8XLv4J5ZVt
kS+BFNtdTuInNQVbXic66YiYb02WIx79pvSPGPbGLIDUEqTt4PRb067MoU4QTYRTjgrhAxCFhxrC
0qUkgjTjSnpBph4lO1JtCH/XkwpHnzw3170wuDq5S/JGrH3YC7JGEgTJ3Z96GBQ//s5Uo9O8uPr+
YaRbOS7nPGvpUea8+TTUbBtUdR9d3hfh2Zl9PsTOE8PhHyxvdFF64DjeT2Q+bjVvH13Z7aH/ILfF
6mmTXksFpA9wbUk9EMkXrUkHv86OXX+8oC5YErkKXXel9XRYiYnIgrlmlCUvP5OM2lFlXQfSZf1W
TWSVHe33ahr6QG1kzTfdA6OWeCsIYRGK8iRiJXIj5smePidbL2szJc32+DaMwcBwfZOU2gHolcrJ
U132258kW+Y4Ac/AmVOcqZOnvmmjQYAjYmZdYobH7MLkN7FQCskoUuCmFQf3WNbIo1gFLFLYCCiY
b8yiStbsRAWZI8skBMKSCdseRGC19+B/RMC+lUtLYb50FMfZDH+LBORaFk1991iSWZafHXUjC9jh
KkScUayG5XxRmZTtNVt0ubsDNL0GY0HhWb91teGrUcfoHhjZwI6ABB96VuFCFihEhdhE2dC9SGI/
NEWWTgT0YVadtOUr20fXXoMUYmeAJbn2oMfqJT5upLDFbbddo8riPqQRAPFsIkoXT/RMXntNygWB
3pnc6AzWbKWWyOmQITerzS/Uab2xqjFNOcjyGk7quzVrWd6902bbQohjb/2bSF6BFml4sS2n0Yti
rYp5rdn57rJLBj7ndwq/Etsm9F3zz7K5oPXzuWSTxBytvFhs85gjItT0WEHG+VnmaTCtBcWeJskU
tRTWLbebBikVEsiFlymsr5dwKY7spm8tsWT+bSkON8YgSsQ3HTgLCzlUbj1smFZro7t5oHpP9QTq
kNT1pSS+UJaOON0Ni4N9MlOKk3f52jp+hqQ0lsP+dqRGBPeM+AQEiWJVmwKBsy4UrL0JZIT5I+zs
U3AvH0eeLWMndZAIv8M58CXAUlSpCQbA9b+rTSyB6F8VfImKbUm0aheNIdypvKLVKeO2zAsLIHm5
gCFcGoep17cky13OIDon+IRF1mR5LgHgPj7YMBwxkDHyxy+8nvkcECLimPY/1R1Urh+ORfg7D8AJ
1psfAH49iMzGWnvB6s2220KgKhhZfHyAqBVt+xCEaOrR9n2NFe0tLxy16qc7wUH1f1iT0C77Su5M
819wRoNf4DhLJTOBhnYWwyBpxBQMR+HBLXdUkrQrFOVm8LZ8fdjbUAfG5xpzhAJvFlO0f9Fl1CIo
CdwlfIe+6uEKgwaSYnfpa1hSMNGJl6jybAp3vabg78yuk7iVaXjomUypQgbWAlTs1cc0R/m4PM7p
ohwLCi76DFCZLIeCDFEGzc8R9Kt9lK7jaEvVFf12iIMXA1XfIWMwawgOyPrIQwv9xyMNB4MMPk9P
cFslfF7n7ZvMrCcP7CnsOWcd0txunuiPsGqcaMn9HmxPEB9yhjNSGmYIRuKajPxfSTas8HwW9pdV
VhTCv3FoEMPBjxsyoX1L8q3Kuubsg+W6e180QwW9VNUW64NPuYWXq0kGynUvpUYQSW2+tNzLyOQJ
UlcdLsibLGh3ezjr0fzT6q6NdY3S600b5EdFx8ga7n+hEVSzPN5HkmQ6ukbL4KcEghZBF8rgj23t
K25n1WQFnVbfe0oCkm/Idl7DX9WzL5lEtzpOVIO5EkTwajcC10wuIFUFBUkpMdulLa7kssoabFkT
wwDUpMwHphecYEahSCCAStg3NiCc98ANdSAFDexxmZZ/Zd6IW7mHdab4wHqySQkAhPnpD9Zf5+kf
No1B3pRIUQ1qD89WF+AG9PeTKO9YlXlwY5+wz9WA4CLF7OIEP7KEOkzFFwsoah8kxK+JTZlGNL+g
a8HkmksscA5gpp6vsLYl/e4lOdI24ttxNRsXoEHL54FyOKdIPPux539N+t6acuBJhRGg5YVHTV9V
PyXwiEv2cMSTI1to1dE+U6uxp0xpBepXls8/xXW6AVLedk6tKZlIrg8t8G7pbC4jpEB+hLIcTA9A
eJAHvcsU//xCgPcDInY7mb1yNxI11D4G/SVfOXj3F3rzIIbzxYKDVK8vgKnVFsWktyVb6Qfplwp0
129F+LvYaHoEO79Ztq928oyZBv3sm8CH3anMoSloa5Oi6Wht3uFczmoVVn9oL6d6/s7Wr5cY1Kw1
gtk/M3nR+50H5FYjtuF5VUqOZaPE8UldWTSfj4OqGiIQyVd5iZflav2i00+dLPBH4xUKpxI6Z36s
MgvlqWq7zGI3Xxc5ScmeS4IoQIiqgTRgoRAFOkvFeYtAdvVZq65vW+pkXlug9AcvwvQzF5KgAf7T
eythfQlXjsB6kXjjaw51g3GGFEiKWlstMEHAeHJfaHaUSTO846DtBIsJWqVj9Ok/f2mrRrTe60b9
TxhZwhfhSVuaK1g2xbXjzelHAjlPBSiS+4PJZRZwwxyEBOdWHj2Wt4wvnRnyOxVT9eC5Pu4x4IoE
OrIKYkT7CNQiMbeaBU332poQqyZ0IYxFaewRSWfj1tMECpxMa3a24B1BGBmQ131eyKQg98xzbbpI
Ca75ECXW8jL8bubZjPirHToD1qyQLKKmluhZvCR9OE2GE+tDvHnJ6zCB5O/Zl89W5woBEt+HnLYe
LuYsQDSM0aW1IdvanJTqWIXvl6KBHTPN+XrAgtmTfcmpVOKrYBYlNadrL0OAmEHYGQvYh0CP44Yt
GJtvaSxaFPJwQxFnLIzBGf4J0pXYtFclVk4sJ2jrLGKHJZfmlA8HqZLCobIxqic/abugCxjJPNw+
0u53diWfdsf1qhzqRLLqxXTqLcnlUr++GGpmngGkmfbYlSunhcl6bbsU5gMC4+bLxEd42Z2Weac3
ivKfv9lWraW+SnLQwUpw/+4JITXR0LaD3OrB6nh/Yyd9S3vW4ZfpBHpAayiXNCcKN/4RJf7vLvPZ
CYtR8eWK3tDY+z0YCADMmd8UecIE4BV3uRo+ENPNuatFTzu/FXwftNI6Cd6hVWeD6Zx3GaT1OHB1
NzyWR6/gp43/srjR/CyFIjNPZJARMYMNBuzGZoPnSd31s+V9sfmosUO8oc6gliDreXUbT7iY4VON
0e1hJz45mq285HtGXu/KFitYT5pR4qxm/4aZGYKSV9sjSyd2BgdZDhkH4b/zYW+xWPmBA8D1H/vl
QBXo7I/AOva19XB/9X4hWEc2/KJXk+aOGLiAI6n0X3KreXnx/xkO8LyCJkHOk4tN2/+VCCYiYR+p
9FOo1Xliada89moIxle9t0P2yarFtdpYMJICJev6xb0C4zvkmJknL0Ag3Hd6WufxvR74EZ5eX5R2
CC2NnhQkhmF2yQ4RXS2+AkNoLn3QY4X4qGwRc43+Sd0URHMqjy7mv5dwvigy/RmhPGGkyGZ/0bgZ
UVXc9xshuw/+TPuCgJedXgME1eYS5sQZLbvKT2bpWw55RnlBfSDy5rTofA2RGXFTfV07RUz9JhgA
bjye97/E5lhgVNexJ1eIohXVqOIVxHUKxtWaJKq1oX5VWJflqIe4pw+Jt4gDDN4plUrOk5zI848G
RwQnCid+TXSA1ktyCyaUiUiV5Crj8iKxaB4d6fReR2g1LZcnk8QjMajgng43dSP8lTgBCh8cdX9U
oDo8wdhbQu0PNe/Px0T/2z8iAJp5bcEvbvI6Fb88Z8XRfesMygIqBwerikzyxC4WK6YhjKFFLL4o
RVVdkaxzkw7kGtLwhrH3kl18W9L+lX3VZevfMhdb3zyMpw4TmmMKBK/dKwoy3aOosxvMcR11HS+x
aq4dwWrp79tNKrl0V6F/kTnG4c0fgNgBWPrYFIVnILuh5SJtONmp+g2ym4jiJN/C0XObnC/+09ST
GMegU5+y2a9yQoPtULAYMEDCpugSA6rbUebusKwDO3PdgzATqWBZf1CyI0WO9AmuqJr5GcOcIbJs
DzR23858O2UsAZ7Ihr4Rq1GGH9a1z/aVH/DLC+Ex5UUFPmcGhC8lkD1aGbPGMweWmIh7SplOfbHN
tP6e+ZfukyoroVNsL4Jau+QolzuImeWNTGrNDcvHTdalv9zp8ePS8Jgq5pKZT9H0Eba9A2XSx2e4
fsFi01u+TJDSyMWoLLSst3K/jtbbN2/YJfW4I8gpbF0bSRoPhpCyWRy7ok6nZxRe3RiXWKtIBNdG
Fo7u+qHKfYTdoy7XrLuVgbTUdRh+iXCWWnW72xQoEGhNo9e/CjVle+tSfLLD/z8ykukvz27LJhv1
XTDIpN9L1avkAfRdm+qXVCmwe0w0roWA7eP40+nHy6siXJBgXNTBXTwXEg6JoCu6GgMCjlQAEKqA
Bq7DwG13qUWKuTX3hPa8ApxoehXatIUTUlNn6zTQKh9syc3KZNcKj7yeGgwQZTXZEzhYJBsnEhhg
7x5neJ9fCCaLeu9LCkGdvzJMTFZXu/Fw+5WHFYuXWBz22Iq/r39F7Cs7X34PMvBLUMEKTyIQcRzP
L7dw9h8bNy1uAYjz90KFz2VrlmIz1VrxLSBWpk/tfyXRc/AZFTsKSed4LLPvb8CXYOCDwfUtFeef
Z2ibaLtf28uVeEoA5HuUJDnKVNg6639rQPF/FtPDh5PXJTb1DO0cUJn5EaNTdf5LbafvPz5Z8oWk
QgCaDdLRES3wBELnMRHv3btIEd/eTnszMrR/9OpkMfPRtNMUFq8RQAmnt2pmF703lf1r9gx1h4D5
Hn307mBM+ReAzlXa+emgaSv1Qsyvf0Ni7QH93IR/P6H3TVHv8qZi0/9QHs1m0nw+U6cH4gDcXmIj
IfBRAIkQE91GVV6Pjp6P/qY74oX0y3NMD6SA0ZP9EDkvqKC3ZGDLm+LG3aomlMvDhdkJV/f3oUBy
jgbZG7c0Q0x9QgH60ymafxwIxZHqsfrjX9/2YntENvOPtbeN71EZ7T/hmC2sUCRsyvQwwYTWqTD0
8/8FrTJRKTfEM3shh7lctpuEBjyc/pYsa3vWfyh/qEF5r3y2CNaafw3wQKW64eGRbwAfvs/d3aeW
ZlkARk2ZzT6PUfcAiBG7ykNxdQB5ox341KSoDJebVwFVcwbM24882Ejx6+zS9RiDzV8NezRHBuU2
r1wc8T+DFlnQ1LylF5SLdq1zCCtw4vOCEQ2Hqy6Niqqn8izX8Kjd7fT+1bquDQXiuyAVVagLDTK+
cXDds6VNrSRwn44A0pVy9YiatS7CTZC5rofBkPJ7tOyGEfcdtSuSn7U2NjI9acCgZKaMuLQjJHIc
aI34fmq9IcskkA/fx1zlHccj4bEA+hmJEYxvJZK96MY3LH5MF8AJNxw6Sy07OKWMB6K7Ba7vIImv
+NZ9NCjbROS4YoeCXQkyoMj00rKx8U7oUqngKbThBLkHRhPxT1gdNAJ0q6Wg5GTyKPMJsPQpVtv+
s2VkQIDqDUVuYXFEz70ElwiRxS9oXUuBetVHF70chRZMDZeV6o3PgXudfIeC4V8PhFG1CmsUVJ4A
O109abd27kPCoMt1+/niWcFTq8cjBNEBhLg3qbJUS3KxZoGs+hr4vtz1bwlRhLHITp7R5q/isjbA
pk30q7DAXFMnLqhjP3yCfn/T+hFzxoRJ38pe5PcJu0oOES2gS9TZx5abGmnoNL50FMpBSefydPll
0Q3bE0qgyiHjGGYtenqy7t5Ksc/O6st+smCACaTkG6zkCl8qDedE1upTE3yDyaV9AvvwSmRzZ4LI
eRTDpVrw4vFC77xUNTpHHyESDVlsW2OWkIMr6AwG4ICtLDAzLtQkRjgqDtv746aYU9zan9+MfnJs
MKHDb+FGbcIx2NlwEPc5xu/l4dhUgNlnIaANxKenornGs+3heAFNt2BmgbjqcZXSGkCpFqhlKWss
oX4qaK9HYVDO0v6mV50UzMOUdd/jwyGWpW7Ucnf+OWCoJ2pvT9yQnU/Q14yH3dIluEVWQ5Tqxz/o
dXq/83j71Db3wMnFB1iMYUoJhZASrTPHf3vHjCPlWg6S2+FLgmHbfBbluqHRLPLX4pyHDwUutm5S
vT16SOkhFu22tfeGhXlTPIqvKZBJ9Qgt6J/ymYUteb0r+iemkJqH4wP4Yet8xu62vpJ5nIoElyQT
wusi/p4PTG5e4lNdDoHbnMwJDjsWS/dFbNAPKU5UDsvEwiqK/qY0RnwOqIDzu6FrFIUULee5YP3g
pDo+ZXZTwZ5UPlUYoBGlodqGdrhmWrdhHVj2pckDNzefvDjbpKZTuMv9xWpAQt2rto7iA0HO6+yc
pyA8pWo87GjZjChFdTanlqBJONUBTZLulcFnJ/hKnG2A2lX3P8c8CSojPDIpats594zzayaOAKIV
f4O3ox2vWU79yydnr0jOczP2UX4TlCbBbms8axwP24l4quSK66THAYWQOiaAU+mJOt3XiZv7zJ6d
ul1P2gQ9gOhAW/jW6hLD51f5vlhIZ7DgwegvDBCMfVWzKbVnvv1Q/YDoDw5CWSypJ2cI+3sKlPrZ
gWdW5a/gVL5jnMWJ5p8LM+OAwOYoWEtT68+ropGb1PTaUkR0/d+FqMRG8ORGRh7EUiye5vnHLcMO
qU5SMoNSTFJVe+xQPJKeGODZAeB5qccwqDngv3yHghHyRtUACB//ti0/sbo0od7bFeMHBzq79j0D
NoVGrC53O0tu9Y/daXvLsRtQ1PYxNWDVucbvdVGNiO/aAyjjoKNK8J/NdvMTHgp1TGltWSm+znDa
1yMYmZIhU4fRAkpAxLFkiGJ9NOzW/CzL4oBKfG31cWEx/K/MLw74rQKXfToEN86S18juRwj6ZdUI
TaW85XBNWEhzQWXgFfGtYlJHlDxRdDqAGjdN2L+zE5jBIv2X6fn00Ci/5AfHieuQG4SkFB+xj05m
Z8kTVht/zU7+JIl/uZD3KWMxOEeGBPp8lXxM0zGvHEhqQ1RCaYkJ6OAetqgB0/TZBFNoIDZ9hmI4
pQoOlqhoRGHpELjlDx5qPg5gZIGtEYi3/iHIT0QeWpYbk5vjm9S5xyO9Xv0uHByKNkPBL6cLfC8J
u6MyLkQ9L5XFV3MCtuIgp1tWORdGCCBGohtiqgxPyUbkp6BkpgoS33D6Rj/0Tobp+he00BaByXg5
EgmMNPQAK7kV6eWqGze59FN9i+9/lowK+iDJZLifNIHEwd9JqzERWxGGB7lRrczKxecBiwI3X6FE
wEJDS4O+MptQ2ivNVLbjcEiSUC5kIr+4qniCCV2TJz8/rh6aVonGiRc9Tj2DEJFwqeJkjoQCjFuX
P2rrhsO0HE+u+KBGXFd+TVKDA5IBrIAEEbjmXH8aRQKiWCp7HZEonzRbJ6I4o7hjyFHXUiv8Kww4
dTGrEXE28lrGpJNMC9dMbAJkfVYycbv0WElPMpiVgz/ARk8iGsqTtR3Uru0/hTeSZMX3amSra/WQ
cAzEt+nXl37jac6J1s2RlxnLsAAUOnDqjuhrKyeJFlqMQ9UstjC1kynomD2NKOpnltY43cHXy8R4
zGV2WRf9b8dZf5su+wnjeoKVUWdZG+ffwkzKQIoI2DjeEZ9jVfsr3iP2u8MQX6w0ivwT2cJ89afR
GRQmsCDVzJvDD6DMizJCAdxPP/5Ku/qurEIXg0BSjoUvdMNdCbv+Jmn8iVFDo3137hrTvIT3HEuI
+jt1H2+M9/nFR/9uF/wa0I2nzJgqLfTjH6Qe7wNuRjO7M6+0CIiQOPp1iBc4Qfzfuh6XaDU6pYDn
cBvXIjALrxFj7homBSsIXyUqnPE/WAtrbM6e7cFL6mOpb2GdKd+O6/DmWsFHJKLC85OvxYJvdaFu
kE3sW1FvBtWb4WyBc3HTscH721x7RGJYO1Z1fwWD+IXVX4o61oUfykzRqnFPXA6xI49VNTz70R8t
+CQRBxPrfKbecDerzxK3Ow1SMDA89TTebujp24RODRxoaxxtSx+U0YsnLc6jAPQIhYJM9NH0eSjA
MYcjfd9SVx5okLDilCUIMzKIJFc6kHUs1KCVQ7JBMkWKlwioMRRocCDYnyW0b7HRbgtzT6Z6USYh
s5N+dwICj7+6uxmik3ty60L5DN3DgAy7h5OrvybZH5NJeOkXf/1/XzBSC13q+Zlm+y/SzfG6nCPB
QwaihyoIB58FkAuN15dLzDtZG+suBwndrgzxi2xFM8/N3xN1kJ9xqMVwOCpMnWYgqb7J4vSQ5cWY
cqCOG29wFdRDNMvs2ap50o/j6PwQOFmuGYJTX3SN4z8n7hEDrO1vHsnYd7ccHWLCS743c8eYNCEK
sEo04GsZ67YF/s0+toSEt7RuN6/gCSVhiFyavKBxWNommBVtSNl8cWjUggzwTMuHYiWvUUvhTwbB
j8GQC7Bh67ZTejdcr0HLXB+ixdMERZXnfQbIEubeCcFbHHtr6QbkNI7hvR+IVJPjh0WHIsbM3dYa
7sfR2oeIQmgR6p2iAXbLptlQZ4TqbOvCVoeRcRdcX3gXLoeFZ3D4yG1uuGXgYrawoFcB8ynW5rqx
3Ci3DRo1kZky9zUc7n0mmaOOBS2VntMjhwz+EWc0585IgDQwAeUlQceXaiVfFGgI/2+xtMdtwTlH
3a6Fz7G1kGBW4+Ipi1UHLfdtaty9WWx2yM2nA3zvk6NOUKqHzO+LK+fBl+B6KeZSkg++eleNHVnW
jspnAQP4Mmm9D3U9UtPe98frqR56uoctxUXc4cVMi+d/TSKPQcBFruG9/8023cUNpD7Sj4WVK9DA
avu4s2P1Gvjio+yDVsm28Hz8rEu2AK/W+xwE/QIWLC/C9o4t0mSeT6qWSCJoWwKk9un0boxM7FPo
13Dxg09EVOXxCDuIE9v0k2+zbG5A2FHP0kjguaopLVXwAXWawkPq9bKA0L1tam2/rY3RdpqcpuEe
856zsLsRGvWW4ywxGVV3NI3RXYZL1pK1YysdgM7oM2qHVBUXWs4y6mwEKsdOtrRn3H9OlGrAhNSq
o0rqQ/JFgGy5zNP01hg+0R4N3TXApfa+Rq7a/66Ds8eF/RLGiTGXRnLfdKEuxW6TEnizY0gQ00gM
mxZgQJRiILJvThW1ssJajACPapb0sk4nSpGC54fp2zdFUK77d20GO1QhGyPki+S6nHhcDQrtecPU
bBBK5WxVylC69RtVs6041tGgvZOu/o4KALps154tw3NtVSXLs+0v+1MxuS3fuxUmn4oM7lss6bzC
Kr5MOLyQUis8EqWUcuw8M9E+JUO5SAT5TdKgz9T31NlFQWPOpzxxX0OQgDNFpat1DBKP3j69nsos
Yb+RIq5/r/a7+uQdzHDtMRGH62Nbis4oMwleYUippWaidfHechCrr9q17QgBtJlDMDbjMIQG/kEM
+9Mro8wCQSgcEGCAvrf1n/eCbGMIRIZRqYjtX43RJOrc6jQbgsuPUidLdxZrUrEHLkEAjwiw4bDK
WZ57imnPUpfHhEQr99WNF5jgWtO0apx7ObDQazXVeDS5jXajGxJ69Ow6TsMbsaPMA7orApig/tAg
m2950p8Kv60BTVqvfqqw0GDsXN3nYH5kS7PbyKPZ4AC4kWmHIfGruGVEzbWfrWySFVZHGpu9qCLC
omLdD1+OygJNlWQ4ubqhHVRH+/JixWPWi5ZaLqJan4z7eVob4pMrBaS69yKNqwiQ/D9A5yQx1SnE
6A3H7/Xahp+nW7hJgnqwb+z4gof39sSJqTHpVoAECp5xKAofpv+RlAZ0/UjIRBtEGUpllcXOov62
dNB5OQEy23Lok8lcKUey1aYQRHOatS+PoQatZBTGBPLQ1QHlyqwx0jm7swcK564QUMsEMRHDQXTw
cGPzAGiZjLt447hc7AoukYWLAVFiK6bP4RPaSUbCk9DpxawwVBv06avrt7gwcE2UZ1g/SmWOz7OR
SgqMmtB65W9ry9fEshHYL5FRM/0nM1ovmSnDJJfcAWXgfWNFVy2eqxhsleG0V+k965N/E2pscXce
fQ3rQKiyA9BORrLp7ugbcR51kLliOye+iVroyUSJeP7bSVa9WhYLQIMbcwL+/HEkiKWinZF5lOYi
tRfxHCe4PdGeeYNrnvU8BLhqeseJEbQlu11sM+sJw1cEliNqFENTz4S84ngIKfWUkaJUEKIPdiFX
5tJlyf8jCqsUYfnxNue0Or/HSTYKuOPZYEKAfJPaZxlVSEtDOawO9glodBUjzbjrVNE7nyU1x/2a
2Rcnyc4erp13OGt4khC3Pi1TPcoi3VgiO6DKxmd2nczMvarRKhAOIUsWOmnH8LeWSiau43QoFPMa
rUQMeBlIuMdpFbkJQctHuDZJxwYflrPlTx/t7rMD0vGtDcJZMEfeCk6mJeTxefeE6+KFfaMDO9Ok
HYiIw+W5nMmsBEtXc26C53VJcck5ygXrwgVp2TMCBlbAvuuoFHDPHrJwoIyV7y2XhaumDm7Vt4vZ
IAqqvUEJjFNsGnm+7DjDx7SuPmShOfyoMH8msmUj+G7fQIId+iUoGXfBhGRJE6kIuxoWLvJlzOmI
qpUFwSniCeHHL5ILt8lbAM+4vo0mmk7tTRHVS+93bdpWTTQKeDhoxpWyBYlVbl3phackGGZPXjAb
xV4YuiFrA2JmxPmGkkr/qRRgLEADS8NFYKOrehhQ/Jsxk2on5wASxAbK/DzIBR75dibewM1TeGK1
Nq/ZHG/xtU3XAWjCDhPyhTa//9g6Z2ljn502FzzALKrND0/v2dR/8SYfV/a+gKtQpiQWVp+yJ/39
DVDfnMXSXYtEeOtGvZPGxLqHyIxXLZwWKnZ/JYQgrrNkcWTVEjbOiZkbMsY8xjJ7Dm/HEl+zQ9r+
mmJUT4Rvq438yMxZ13bA54DH9hqQQIl0g510GyjU0F9qKdx71Jjo1QBJkp+HJMXouKyh12KqmZel
kVODVwMHhnyfmZkY4T+mBkb4n8of7GE0S4pWzYY/6pWvgzSsKHoo4h5zl/3MWNsMslhK7Xsoxwzs
CZwKeHltW8r0duE7H+kflP1E7AbjauORz9QZ4Kkhq94yjltPPvAC2M00lTRIxUrFHBHUg5/VOMW5
1aTYLtvRdTgQrL62mUWtIz7fx6oxlVSA7XHGe0hzGzAbybRiKL7rAmsKLa6LY32Foa3ZLKD0byvN
e8LmR0aFvWGOnQ80k00/FQrzskyo4KkjDL3SUjPCn4kNYqASNch8D78oBCo7iyCV4G4KPeTg9xD6
rXjSj2qTn0iLKJfdYApVIO1ZsQofsMogYDHWVig4NzMe0ZXbdWXWRDJwllvb9aIIHPEfajGvFVOp
WTH0OcwwvnwT0g13AZly2IxvDRA+4HpllHztgr+l9mwOVjb9CrskSHmzn2qQJgWhoclqL5jGSH06
gZz22i3WPPembZb25N/wMZ+Nv9OdbHJhOB1rHwNyatKKrSkttXq6Fks9DP1NbUoczgkHnsx/kcn0
HGsyNVdtKAq3/Zy1Qcq2gbEEvBUH5J7dTFHw2QFifTPCVdBF1kkXObDXF1gsSUsI8xfSjUaWumFX
dsivzbJZrvmvYiP0OAordSkkC95auppKDROOcaWTB+ioYIBTz9HVZ7HhzBgTKFEtCNghKDlvhWFj
BaWjIlmdByReUHbMxXPseDihh4R7kdb8od3Tdyg1H7eV8i8g0WzfXqNeM0N4PQ2kl/MAXd+8pPki
yMPThytP353CmrfMrvC+xpJnoNGGZfQ5IBcSTrK2AOZVUnJXUCgl/P7Y4RTROwhEcDLiQtRKfDq7
KyjC5sDlxvc7+b7gluZ9Ofx+D8yJn2rvo+D49AZGF2skAX2ktS95mLMzWNlzKhNfttKXpV5j0JJk
HUlcTbYM1RkCCtu5yepksMiosQtLCHhR/m4zMFQm2taiRNDyP/ypT1OTXJyO/1j5zXOp6YCm9WPf
wgn6D83LCP39410V0cYDi1hYy+a/nzw7nTIsOBmhDvPqAjEl5RDYFZoBEbPXxSDujMNp/guoUPfD
hzfmPOuPkZRKhZhqAMQZy1y3BXurbftmijvMN8yx1BwmmC8h5jL52lDQGfG6i2EMfZqwYUksW/+E
MFgf+y2R+tBMydwQYyQ2pzSIpE55AQ/zkPMleF5k7o1SaAMSAccUSI3V+JjS+dEg1LavDI9k8gOj
yla+im2Fg6URHfRCdOl63ItscyYZbA35dE+frB42Bo9SEhm2opRnWzlettgz19KCp4S1fHCcoBi6
motS3pToHEomh/Dfr9VjjHqU9eWP/frCLf7A2uZxjuTNNdm28wCdF3256qBuZnqItiL/sz1WnvTZ
3ps/GfTP2ZNo1c/3jm09+y4nLH9+udaw5pNSeyfulA550U6ppxQ1Nx5/SOlMfPYDYFuIXoZaSxRv
PSv3jCMFH5bL9HhtyQzw1E3o5a3OqeBiERSovE7B638r2hrsj5O+iW/zyy/kiDbYSmGiPMpAAf0r
hjAtBIlH2/N9UkdoeDr10ohIMOiCZ2elgu5Cf9Wqr3ESzick9K5egoKnkOltKHDT3pU3wnEf0XSZ
uz7sv1/mMfCnEcOcOoBATMH4SGk+wyRo+eww0+QCd8XilKGZ3AK2umiDip1j6+iuuDx82mT9cNnz
ZkvPB2JcCHinGQRX3hRzgZw7ROYZauEcUBvBcSvlR5j23sEhySO5T89P3kIjoRQVnR6Jkoia1ZHD
HltT1vqOCX3A5AzrRtdQ/KAZVO+knbrkNru+xvnVZ8HBgy+eqipokhIZQO8N7gcZnSriTDW2/g2H
AQyJnZ5ZU/K8GqUPC2vwm6oCzFSk7K8Bwlvrz483tTU9zEMK/nlr6PWqeNKu2HlcpUOy04BbAI32
by7i3Gj7VyljAEyK+zRiQrJ4Aox8LxbKcB8gJXaGZtwNF646kYAe+6uM/B6lVQ0k3GCiRZOgsvst
84qRY2GcjfziS0TBuhB4baRwyerQzAY5sgVo6dPy8zMyeMAkFYcGY+ZA0VT4WqdVT5TOEy9sCLkn
Fwuti3cPhj3fAC/AYFfdq9ePaw4g+FlzIeYMrh64l0+kxS9oY3FhlkZKBZcLuEF5aFdkhsPlLgEU
7NQF97HykeFllCnuN2miqkIrh37E+0DWU1ppssxpUmSpKoN1poop/aJvxPT8S+wQoM5xLXsKNbR8
0q8ecm/lCGp5bOZUoHxoOp02c+wDM8mZWynwZHIoerCwZBi3dq2IIF7luDTu+dLjN0hl4rvPVSpt
zY4ET4PuaR4ZIqsJPhcF2TePHYQTWqsFWtByCGxr+Zdu8bw2wkDeCpz0REixvE4+WPFc4g1AZz6x
OmXqI+iveF6R/LFfkCqmZzy5hufnCawrxwpCQ6l77riIbU3i/P185YDmw75h4gaX79kUAB9KFx51
LGUO1Ezw2Mg3u4ExoC0Yd8KhjFBm/ca4MDPOqGkGO4f0V/ZxQEmoZFr+EBS39/juZQ25IMJprETR
L6JOFiIakUtWF5etZr5I1X/d1dF3lvvUJysXAZSqFbHpBoc+KWy7MpbolOJaTLsnItldd0Mkuk8U
mrBvMsuifSaTySyN2jf/Aj9H8hzAB+aaxHfihHiZjBBhGNBGgMsY/6vvTTGZkuBly4VCIBg0OSdr
uG5brhFiLxKmqyZzPEOybcON9vFr3GFiMfFLkncBNNqsyxbqxE9Ky2ri8NdzXkSO+1+7grwhQaxP
IoQ5rxfELvB69Df35cNoocFWhWhYIz+HpSZhhLl+VyRlyhcaooS8AnkFlLqrRa78T/4j1A6F16pG
74RerT1J0kEz5CimnMaB2onpUhrVjE+WLye6ncPDxevlPxAlAkz9tFsQbPiaTrdnQWWe/J23wg1b
AX9czSdU2DV22Q3bny1jVCszg9l/dyda1V4Ywf8QmBb+Wx6UWGYlxezH+WCDTHiRnoZpn41E+bjc
pYSjvAMvOyRMSIKDRivYmwDazeSSB3BCciQb+2mxcpBhyBH4NsmzhvWC+TRja23++chZt313Ng+A
wVLSdOL7mslUxWSR4eilGob+P+ivhpcMd9amoLtkOQU8GBBAnSodCKRwHFbsT/SBDsED4WSNyHZZ
Rtn8Can1mEVu035BlM9T5U6sndRhJTr56KCSRNKDM/kIdP+qDyvu0KNMl86B9jumNc9AYe7Pe6aQ
FsLK9NkWwiekN7LdI1/u8M/o9A49Pg08x+j+Oam2pWooMrX9tXe9EULS7RT2WjMicGnsPKTggRaT
aGsCP9ZLeqzCfnmOuYJs82hdA3LRdZfFE/U+W/b1ThQieiRki4uz7mr/VvT8E3ehpONE9XBDXMfQ
42dBGsaDubOtV7+uh6WFF6OlOAX8uiNT9nT/vPxEiC+c6S4iBhMZoS0m+Tk0BA7nIX2ObMoauk/b
gB52HgNW7GrTEbdp2nMjIh6GMU4M6viYNiiacq5KJfhHhidV6UJiZ9GAjlZgMvSzjLmcZJJlgTjd
rPwHvAQQSCAwKBHnCME5SsT3xc2AQ51GW1BXUKQls37iP3j9t624XjcMQkRrF5pKQtKe/h1C8hju
Fp6VqE+v8Rhh3GHOc7SkDKoYzBRU4XlnKgKlUMEzg5y7DVxxBt9hisa+S8lLlVkbkPpkYlySuQJN
QK4ztVBNKHUzZCmSxYtRkIASTa2sv6j4iQmXdESufYoicw6UzEZy/vJbZoiZpS5ePEY4pRtTpYoM
bVt7J4ZmjNx0bXEnEbKwHXlW3PvWGbwkc+RuIRSe6GXwmjqQExxAfAUIOCxhYr+FyLydHsWLJMNp
oIdHvgP5DSoO/T27MFulL8XxSk7akVgr3Cj9S2hCVLop74ZS3zFjgb+xfVOy9O8a6ECA26PU0udu
uadUbyyTaioHGomo+d94RI/0SiGG1eIU2l8KHDBMYYej2JwyFrIGBMJwbITt7z2aIzh0osYcL7CP
WqqFfoKsRgBykTG+tRI1lw6oKKFhPg40hWlKgJQEJGxK57oseDPeP7CALPQS2y3ENZU9CzyQof2u
XihzVgAaU4xMgnU/NIMqiHSizlO1Y9et8hcaUuQJ/sU96UlOtOIdepgshgRay4E2Drpne8gnW7ha
H04Q042tHHO2sEc7vuYwe4IOuy8/1xWyWhOXl3Q2vDKZTZJwGv77agLj3seg6Gv0A1NQGFG0JS+H
tfU7qLgSU5QjZVom6KYr8YdtHUktaSUyw4daCVW8qv3DjKU0orEu7XMBgm0QdDllV1n/wCEGs/Aa
3GjX4HFrbHjffnD3LzvJnjlWtmirLQNtzx9+fUcNDfFGGiWS0+6FH2RXoJ2bUBFyX9ZFNQcYRExi
oRwIm6ZS0aKsff+3R6oY97kpMyh1geVMzJGvy1Gp4q7hpYKMDj2OHLMFsKa7suXct4OlTX7edJFc
mQvoLoUFGxNseIcy6q2b9B8crAyXdxNw95p4I1ae+LNvVhxBsUbXXOzkze8bsb1fGJK9yu1DxXNg
EGeRRPg0g7aUZNfVkxEM9hQ1aBaxylmAna0P/31PoxBOel41Tc7AlYGbm+DlscNkgdo0XF4L6tdJ
9RYtLhB+l+CilqeVml/9wMSuuSTHHg0jNoknxGOQXJhLf3fuNNVI5lUA5A+tzsD3fbEgNjnuZ2Ad
A9sJBnEe357dl9UbJg6AzTBFKnppI1O0XEtAprO1/gouRcDZrZh1FqPyLEwc0RXC1Ojcf3KnCiY9
K3g6+Puaa8YnAHSiSMref1sAjx95o5rey4qN+6ihELMk8/qlmqguL+lOEr0A9a6h1BSyMrDTiPmp
p1C+Vk8dTqX0XF/mxjYibvHB8czYt/+E3H8WlH9gyeICOgL/r+DgaLhrTtyeQw0soOdDsBcr7YTG
W0ZQ7faaPs7Zk3sC9WyzjWAJ/yG8CcwTxTdDDKQWW54YakmQD0Szr9XMy9jsn4mXiC5sbZgBk1cb
Ld+/yw+bo95HK6VkvE6lQQPi/QQnJiOqCNQLgRq5sVUqM04ytWM+pk3wZBHx5oVIffGJgjVdpjob
vdAJdjdnVMs2yw/lXWM066vGEaz+wOubEnNtNFNlSEmI7oJofttWpsLBatXQzanroXX6FtrCuPRT
v34rD0CGnu2cJSwiFQMZVx6I0ED+Q2H8r/JIRs9b3ZHlBWyVs10JmmfPh4UkmSDOHbaFRmFqcXhE
LAjEqAoiwdVRC8YD1BAv1RFfb7543VURSvV1mRSV2SaxMuP4aCRwDiZah01eYjVXc7aqfCYSOMF5
ElzTo0shHleYOqueI7j7JmdBsyrA52rsZeMViN0jNv3SZ86KE57ewUW7MvD5J9J+vz+tvntAVmJ3
FO4M+ISxvI92aPyEQrAceUtAIEfBL8c8ciHe12OHY32h4G9JFbAGmFfGloVJjT9xnd1qi+kDZR1c
H1qjCVbDBVXWzp5BNHNMMEADwFqNHCcL1nYuA61QA+FBJ1OjShXUvZWDBsnf6sk5LyVdQ6Pll4fW
n/wOgqkhBdMHLUh3piKNeoR81FlFVm6azFPGZyZ6ZuGy5pIEvH/H/ruTy/vAwvdddEeUL/+B3uaS
yE0lXgzyhADtDFMRlHHlImWbQajbHOtB+k40yMwovx5qpvdQx+0FX+oIibL3VuAegYba9UW6qPwe
hv44JgmU1qFwOsFu+6t96kYV1mr4sfOBi5wr9Z6emZOR58Qvrc0sc7xLp9wPg14c+vsLzJ5frvGJ
ks1REJg2KwJPOvw73G5fNABk7WKc+eoErGsy8lT6U3IvZTkxmxP3IJvolziJfyVS4Stlz6jxQTvn
b2+6KayZ39OlmK+LMphYVlEq8wyhnuQC8S9EiWnsdLmzP/IBnB0YYazt1xPXwLXCzb2wK3OUIGIb
mHfE7yve/sPhMvDB8Z3W4d+y6FpQ3cZJIYqc1yXtlDR+ZagbR9kIh4C3uxETkLrDLTL26GVEpc0n
I7XC7cEQEpuZKHcq/gV5lGIEJVODaKu47Hd5o73PvyD2VoAh7ALFtn1K/w5lCV9nmadzOPF44yBk
Zqg4wdUVp6MhohS5GcHzqmauWr9C+10TgX91h0ls5AT34ayhXUsqNYuwwKlkSJ0Cxuy05PHfp5pd
eHxJ2edq4ExcZ6/YIt1hipqCPZsbJu30PCYxOnO+2Yk+tsJNh9IIpZ3l5AJ5BOJXHJkiDpheZULY
akqpAO3dy6vuysYt/Gr453PEqoQlIae4CugueC+doZnzX6v1Ig/D4fuND71aiR/mDFSuOjrBCyVy
8TMvZKOKXUmLfkQdUvGhnhC7nxDvTHetdpojo7GLod8B723S9+4GCHtQm3mj9LYOTpjeiQFzhCwT
2melX0XR5YBKu7CYYDAXqCFPayugJzzn1J2XJEMpQRUMimxfUeMiQb6jNUUSrrFpctc7VzSgSP50
ON5eBt+evuTS+VhCqHsWSKGY0+Nei0pBWIn42rK41Prl/iR6/lKKHj2fv7SLUsXktpdVgrmic2Yt
5VmujuIHiiGqrpvVFn4nLlND9yQJYmAkQnoSjkqQdSDusw69c93PEECcjYX5UBKypWh9MvKq1VGc
7inqLRA8nKeb1E6T77N5zmcXdwy4sRx6L+QLo+OfzjbYbokEPfOuPRbjPvZR3/xshXzaNddYtfvu
3owKO7isAVfFfJ+rDxwNw3Wyxx9ZGD1ZhwwbgzAMRJj13sZuWFty+otyi28fizL9aMNpJsqeed6G
mvGjfWFCs7tAq5eQiXT0HAOi0Tx2hEdUXWCvyayrcwIxQGBnmDG75kzFvALG0+MuIxt5IsisOiKd
X4eaM6N1cH9f3CqeDB+J1gEIDUU7KGbnYs4aXDE2IovvSvTsoPJVJXrpl2fcLwIvu5IwIiHxZ8tM
4l5nV1nC1t72W8vRy2oq7/NroflJOA4iNKBgnbcO2tseFh+GVi73vSZa0XqOzlqrO6n0I2c1ZSuc
eC1xqnUA6HO2QKSH2E7izKI3USmEJY75Voi2sPZBfgWNFfr1UhiOiqPjcM4ns4ZOTEOJdIA50DZ5
H9Qk7YmJlSyE4PDPlrm469k9gMoLYDeMw1JK5oVnv3J5god/ADp0TVmPRAJQSKE4jIz91sK+vXaP
nl7L1PPMnlQ89Kz5HDHTKn1/SMVLBDeKXGQWCrvzcqnaHuWuOFTr5URb9dHBha8QbTTIJQzlp6ue
1ssD4q4fBDPMykGszR1n1g2AS6dIU9rPVYXznuJCxPLF2BmjWhzvoyjwzWhk3ORndLP3lLfjJiuY
h4OVp3BDbQdlAUYVtmbHi3bqLOQQYep3CvwHqt3yUaf86OJPO11i22PUjpcXHfVz2PXBnyeDT5eI
QS+f48eDCKiuAn+UuRMTy5zeb0CjDdjcLUqH+QJMvVhx98JHg0G7I+X2kTaKz/fBALrPykHivMrG
RgK99X93/6AMpbVh6/LjEYueNefGjnSozgpsz/dKAwKFzKf+DMfIrlJuKwyh98XgCxv2x91V4AMp
oLxhI13AdXxxDLz6HZdFvd8GcA0Q9FzErsa9jqjvhd5poTR3ZVsgpliNEdUENbYaRQsjW716BrVK
4gKXrmVLxrTxzfUBdlhjsFSzcs+QRVUOTy1hL0k0/r124aojZHu2W0Rq8TUSCH1taDtzdt9HRVDL
qJHZ6ZOo7J8rEdXhW2z3S/XMRqVxVG0KPR7RkHKhyfZfyhAV+WoyTihm6nLJWs+rzGiPeCvmHTFG
L4bRZU20QK3MpzOVIpmFUM89AZ+JGzVgyY/kp5yxBJoJqjXz78tnqUR0YmuOiiI74Q1HHgIRfleA
pkNn48V0hEQQBzvlC06HdbBkrtO0rlwhTXR9ObSYZO0QzC2MbKBLTLNwDyMeQzbIloxZnBOek+5d
5GkvlJ5pvnc7D91aHLsXmfv0MbnzzYWJxjUN3tHNYgXUrAOQhPWvFgEOTZSAMtaC8NtWBvZVZluo
l0xyNAJeCKy8nYWdMVnl2Iiu8skoiRJwZzTv/5tAStxA21BfocpBgbMbSLvH8Blb4aJmja80UKX5
ErJ0jWtYlmmxzcKJ5ChOsFjhA0yyn7JebQpWD9XKIoonPTckTMuiqMPEWCxCd8AqnAptu/FkMsGw
vdipjLCvTX7B6u2eyx8J5/hEAMGgl8O4syyf3UzIALfQVB9VvXdUybrM5ClBabccZD5ZDedwH9hQ
udom96K3pjMECLbRCqk1Zpyp+J2dI9l+p053+8pjfrvG8j2SIXpuYPZA5g6H6/Kl/kom9XFHdj6j
jPf724TaHO99eK20WQ3S+a63ZKWZ0c33pdL0cBsB/rUlIFpnvlSS59BP6XpI9AGETEOBHfRXjrd3
oAG71UUwa1dLbrBFs/FNEqbcDeM0e91nMHC+IgGdu8XK0A9BlfocwaTZjh0rzAR+o2pvZrGEcz/b
JSDMME9O+TZeTXV2NVoLukffeNlxwkc1C+Qqp+CkvNfVuAVnrR32QfMf6/7+yd7A0EvmuVdW4EXm
4AF24El9w/UX3o1I4ePWfa/x5ZlUyO5kT+Lv44eNISPAIG71Y2bwk0Z3GsL/X9DSFKJxXuxVTVUl
f90+eqnwd+FgRDFvp/B1g/hDfc3NrM0A2FivrZ1lVqSWA33SjY7J5y49UE7FIsePLYt42LlEE2xZ
Ud2OH58rtBrPtMM6WElOj9wxxltWbCUANH028Kouf2ngBBzyffHVw353IfVcqoTVbF+768mEsDIs
vJJWEWCoLER7+C4NVZr2SfyDopH9nuIF8JgcaWDJAjcu4+6R9I5lcTbepvmkNVKlCa7Y7/aMja5o
kyFStBqdX76PiXe0HIbomhzR8bWRUfpWQFD8By1dGtC7qrM+Iou4/mhvIpFWdTBTAhpOKwH1YsiA
8y7OP3kbG/P1H7IrnBlzKEAXfpPjK/Y0B50smkPFBBuV2aP4HedK7KERSXKyGwiwoLNOXfoyLE8+
s2qWKyKD/bnfGL5+esv+81c/IMelkmOBle6n4BFuRLvgdxnk9dpmyANlSzC5PcqKpcnf55Tx5Tss
IZIQZIohQCX+UOvsJT+6atNF04+LxhlNyNUsacuiAdq8siJfprZTtmid7wDpVVj5vEU4ccJx021v
AIBEjlglctRlD3Z0wnu2qhwzYpza8Z+goZfve5bktj74V/+z8wTiTG5VroyPb8z2s3P5zJt31rxk
oIiGVp0S/TSfAR2iayc3403v7H0A6+2FCr559iqkeF5PD7IfogtI6JCtGaGsS2VZ5WVo530fvs+n
KFGUG3KYsj9gkbyHq6gIixuIEyOoxhBompAoJz4nJhBBO2mfLqrDohJb+C7MOY5Kc42yvvvIx5Gz
s3zpX1TTLaiHJsxERZ+MTXtvar5KbAfH+arVNej76LMX1DT/4PHBXiyxy2Sy/hhFZ7W1wePXpDlu
Es7ZaR6c/5oKReq+pF1A5kSR/13L6MZi9YpVVPcZMzdnDKF+mbxO2oGtrSSUsXDcPyyL0ZCa361C
54KoK93WeAnQmM0QVsi3bvha6gY4glqWNmDgQzCZR8/194w1ROj+b35Xaqy922Ad0i58ixWJ5cB5
rR+j0GRSUe4VmPwpTltImzWwHpyjNZ9TTd0YnfkZGZ7ZthDAy8DXbNBd4JFQU9p9eAzGP/QA5qbr
ZcUipkf7XISJr+clflHaAe5Uhu2a+l+Q2Fxvdjg/pYNgbnoR8PmAUWrdtB64AkJf7Mi+NaDwpNNb
LEZq4O0fRi1QAe2IWRzayvhcJN9g1ox9oTMzKq0cEe58kW9qbK8l6O8pSkcMQsMbP/OPVeZcnBqZ
kFXKmrCXhN84HFkakZQTId1IKHZ2IlpRtmv7mR/UHfZ6+eHjxGwi47S7oD46+22tHXXZMafZaUeI
eGZkkQ+r7BOCi66/9pui1yj5pwZI9p/6oTul3hD8RmQiq6gjU8g4hZgXn4h86f5d0W8mI32+PFNG
ookrmfTaa6CZZQw9Up/jNsq8QtMLJnIYIVaB4m3GxADnUNdoWpJKY8cPhs32hIQsuhINGqipPlAS
fTBxBaNtsBI8bFp8tnv3FoPlZahWOhJgxgHQa9TMzuu9OLMQFtPfLee9hvJ3kFiao1C5h73BVNDl
FcJGZpIGrz3btRYhUYTVv9ukzDgs3EVF4nStgGAXJ31laICo5s/MukECi8Ps9dcgWy6W8j5SJ0yz
dHFlO8NJ+d/0VJn54fKx77vpvmRBhx3nDvFaAW3d9AUXkHhdcCQjIme9Gsl6f2QfAsxNVGXeMwUG
Cc4bTX4m3S5HBxYnarLO1OaMmxT6A/1ukLVmBhdUREDLsntabP06M3PISoTcN3UcxNuUhUf5BSUT
eHHTCzrD3QMAA1FA7TGPIond8w/DiGA9LvuPSWtnq/0CiFbq9BKYoI7cDXlfSFBQtvhp+gEM+FTs
qiE3GYhfedKUwHuIX/sG5gXcKVeTyhlW1ayV83x+am99SHNZbcOqjBPcsjg+OolUOgolbo8IjD7r
9IP1W0gwuV8zqT3A0O5fKST6tmyuIXnfyqRWT/71QFB1o2tIiQY5Z1HLkJYyOPqVfBbgd2bE6izz
vKyfqW19BVa7eAmxJrQIlX1+odfnnUJ6jgYnvzikssQYsBiKo+mUsFySnYM9RwGAxvJqGvuUHlpn
3vRpk2BtYOrxzRlt9UtMmF5GEYamckyk8qelJmLSQmYd5zZV4PenUK7NSZOQxe06SPUYQq5d0iIU
AjRajvzUbou3hDCW03AVjr2S7+1XY1c9Xub1yAsds9cCbxndGvnTzlNafll+PvaxigxOsspIZqjf
4aqKxcrPM0j0SHwopo1ibMXavrSq0lOEvoEbplbeWDABY/q1gRaRVw5EGD6shqby8jKiLXlCXcMJ
z4v/CdeQN3E+au/a4EqA6DN8j2nC9Jn6aNotXvnYRVH0JBdTyeNjM9A/EvlblkLw/XFlaLWmte3e
pudUWaNPRT6naoX2pYblUu+2aB2V+M5J96JpyyPRKMF/4tia4ATiWAKmHTkvX1uOC+9BV/9lqilN
lE9r785M2v3GROXJEUdg9RCCeBaaecJ4xe13CG3Oo1aEsfpwQALHkm5F0ExBHV2dlytqVRdiu52H
Nrocn1fh0zR4zNVQbXTdJ6DmkcrcaqX6wPGjb4W3EjSYWBfuOeBRvhqVuR/WhdwwoKSyHahup1Ld
TdIGyjS8VGlJF1rphJgnVolchMvvzEmvpBCGnRWpfbGCpYb7PPI4PM4H6DNLF7JGPPh8Gxw+1SYH
PaUfQPAG/qyyLmgsOSShvTtQQE7R0S4aIGch3H8sGJmJINGLddT/GTvLCWTna5b8iioSRgQOSLLj
7voi3PlRq+MMSqmyF592SwpOZXo60JYf8aw3cwklY88W89jdipvu+NsvutIWwH0nwOqaWNtpfSwk
HqPqTWo0nabNuvnf8z5uattlwDw/o3pb1GPk64c+MmZT/Y+QfztI06OuuHdAvJI+9FeM7NF4v+yz
IEWSkEFlPZLzGyMfISleiIDCKicngUeQbmWFpYZwyKq42/hUytDFjgKIybGqMeodYLi0SCRdju96
mS1AzQLJrmkcA8LACHRJkvqzMKD/5swrHdLOybo4OlWJ9OHoaEy9W6j/+HJJ12aVRgNGWI0RvW7c
tOJRbHAdtT3jRP5pYwdJUT0t3q6mFnLxlNV+c1odzlIIAl96P66I7cTczveHlcRhf4Q2PVezBYHl
ic5ynUzAHW63nij+xXmX5X7Ct+fCuuY2puoQL/uYU4pAkfQbBxJ1eWap3e1h9+8BUIlkMlYZsz63
cFIuq+q1TG2H7EvejJ//8yX5Blhjh6aVVxvDKCwP4Cre99cEn07wOTgJEKBa6SZtqVBxHiYSieEO
z/dYqYHR06A/TIUw9a8ULN2e6Zy9/2n8D+HgwFoudjyBj83ie3MeexPXT9nyCHstioCRi1HMMPtb
XiIhDIr4v0BJmE7ClulLq6hrWDoRerG2jZ14xxp5BWSJmt+YUAotCpbXSYIJhSd0myXdJJOB15L4
1dv3RL7oXVoyCoVNkIfzcVv9uy8HVlzgLUag+8L5WvAUnEl0Vwf+ny774YNLzw5+zoFUEmZtQVik
1aCn/PtKII23Tk3qTKN/YEmPmp7l9MP9Q/p4wl8nkOgpfurVChxWmVtA2CBoqa/LJV1is+RjsoSo
3LZCyAQunMIeGbP5H4HjKSwE//91V4mpV+egbrTgcb78l6SlqA6Gdcwkk/7RG/SuLb7xDNKDeyU6
4NhBjdK3LYTBSp8DYY3XMQeL9ZQI/4SO2FozUBB16b2PyNp8tK1hDrF4IO8Qk1JWp3YdkWYjI0YT
W6a0TvGic2ZEeJiI7D/PGQUJjs0YNjWc6lpXLcnrDRQkC6nx2hFTLNPt0AfDNfTCxEDm2JPgnUW5
so0p+iZYiWd4nfLORJHoLo8AORhJOYocddAR8yQP64hcFSNRIHMQqg+Z8bZu1TipmpGkEVRhcehd
Klfy9BvkBHDO//kLb5lEX89t369IkfXgpmJMVxcbUtz/zdlX5oEtHwnGNzxm6m/CUg0C94YkyTYE
X6T1PHwCesebgY/91YagoFOPVor4ApnvHQQVl+NjWbWjF2eiPMd61Btipr5eOXy9qeKBPGbuVIAN
nCR0uXtEFa3eSWka3oreew4P5RgrzM/2O4Ee6A4wXCzqPbySZQ7trte97Fv1Bu/ikd9ymBuGDjZ4
/hUMf0CGJxqQpMhk23pEMbAfqT8dfL2/vcwhHQUpeYFHtc7UiKhmoS9GA27x84eyxSTR53GQHriK
18bpmWAoJM23XxLlW5ZmGK18pwFOKhum0QbO/ecVUAgY+n2VLnn2P6NB/d6VfIYF079I7VO05UvP
CpF1zVGqu7aj3kDWtifROeNJ8hmur1nvuWMM7+3OD1DBf+f6oMqEWISICBZOpPIWf6Ghd3VJcYZn
qEMuThcgx+35Q/kLpm1dAoZPGmcEGUD3D2DIgqwFpj4TQpx+csI9/y9zH47zxcP9ZksFmomKVP0r
pNX3l3BFL5VNdKxuaH2JMRYDRLg3J3+38h2AsUawK1T8ys5M6Ae+fL640mZ/ea9VlHjHlTZWTkBJ
aXbR2nmSouwFr0jtxWohe8ZOxQDr8wcA9MyRbURAY+YG4Zj110eR1q5gDCt9afA23qYJOk6xJOvK
sE7OwWbBPoQBCQhHlcJLmf6PFr8kMAS9L198sB6fstiT9snLJRCf7YInR7izt4zw8ipf3avIKYpr
gIcrmTw9moLCcsHAQmAojrpKlDF3CIv0K1bXJ/Yk0J1q1c8D5XmRB9b85PZ/IfjkGtOeEcpI5JYD
Mzy2WeepNydRuqsjW6JmNhlBolG1krakzUg+DmH21JmMzpmnCN8SN74tqY9SQapFqhvxZiJFvhak
dSCHIF6VkqEduwU16wz0OHXz9jpeBxV74Cgc/pGyxYsNgAOTjVsqDUgbfvs9gwsAhD0e7eFiEdpu
dgiinT610cKhseK7D5d/UaYgIGOnqS2IT9vI13V7VysP3GHMDfN8FA70QvCu4EVczhCkiDvLxrJQ
GypRQZyAEpLg26oTy/M7egEnOzAk0Jq3SfbOJrwRcZuTjRh/3htu8Ks9s6Ao7kZTyttjr9KfMYFh
M+fADD6qzsEeKP+F1el6DL2pVE6XTLMlSxvxxst8tfUiC2z6lcz+DBXFenTHGikcyUXekffjjJlv
OO7j6SAoK8RlaEY5/XW9uAXXIyGa6w59j6NEnM30jrpp1aB/olit09YKy2hZmMbk332Zy0yeilQ3
4vSVJ/oS7mc5sxj+nVib5J4iHwoRsRASvDjHjo2utRDpoEN9IKmjxR2i6TCGMkZyOSXQ01hO8Z1q
DAk/NrNCtnpUAr1SJIYNwXp/vKaFkbrOwm+7IOhFpe8XRKaVI/ULMpZOWvHWY//WtWU77fjKfyUL
c86Vj+xc4cT+fvVf+KuTCqcR7558/O6EZFbV0D3zOxESjCJvBVkpSrnKTnewGswkM/NCAg3ve7rG
Hv6Lk60pLBVIEmtsxrQZGgROly7iCJKKptTCzQx6zLe4bZkuPu9GHDzDtb4PBTGM/j04XmGjl7s/
w7r3t0pRENu2BfnkFXHAuGnP2C5lFVkJi0SGLMFlr18D/oZ1WcMT/+2qsnH6HGLY3fBUXioiHZmj
IX1uOPMe6VhATomkKuWTREfd/2pc4Rfa/hHdBk/Hc0JtbsF6mz7jf4K5p/OAckxAopUzWXf/b6Fz
XURT3m5mkqebban7WlbtYeYbCOuDNZ4XYVB/CfXS9Pk+Glrb6OJF3L7K8vwKhW5kqo208mWv/TRe
b1MqjObUR3L1RFiMZRkb4jOiLBk1abIwQOBcjfnA/gnOOEF1lsje3kwxIV73DhLPoM3cHh7HHR38
FbgyZE1dmjiPybXdfopCxru60wFUu/TRfa5tOuAuqrSmO48xjirA9UiZEyH8MyJ0Ortg58Y5S5yu
YzTRsjK1ANWXW+aSCsGqBoh8wPmtJszu0hp9Bdvd9sDObSqIjIBnSr4qbkqPOTs2/3o1dvQg25Nq
sYS9ZK56x0aI2EC5tVc33ERWawNuVEvILM+LAnLIBayMUc0uuKe+C5WzK/7Olr+QkpqxdKGsmgCL
9o3Z2ZqhMqrJFdWEv5h2cK+bL20hmkYWQ75gq1WhVk8iUXxqe80vjX6bfzIj3QXgtWW8Bw8dl1hU
t2d8C09nF79BvDIEqwp4A+aZBOIuqdShb3bvrZytI2+TiyeFuJGjM8IX2lntX1As02zXulA0x5Y5
E40iBri9cmtVKAcTGC3FFyF24S9t2woOLYfD/pqs3qHiDIJfVTcFODYOT9Ry5k5CndhBPOn41ro4
7gYMx+TcnFD4ip90QQDsNurlwioCbI8CoSrTDI8e3AqNMT8JGCirqbVEGL/Rw6I0guZ3rOkzhEAw
a92D2nrDGFRnn9+mDaREJjUgKkBjXsQ20GvcbrJzl/KndVhteC6fvIWfFqJ3llEnoGjbhUNi5k9I
ge9G8ihKTChdVls1V3bZFOOdc02qErNF80c+dH3Gjve+NXnfWIOa5ZYj2FYW3O3JklgzeCRdZsJF
t2FtDbEiw9MRkefHZ4t16ffJcmAzRGKHIyN68bjyzZHxjgfejChyz3ZjZjeco2RqHt4qU0sluaET
FN3Q9/MpGWCIqHh80iodoPwEIN7K5kE+mCsaSiyA4Gl7ONo4KU0jpnHYvu6WJU8TwC80KO0pXPMh
Cg+g5ZaoE2Pk//weRjuI9H6IqPtpm0sYMydsodNK3eOOH1c3eaKYDmai8IK4fH2B9yr02HZMWO1j
eZ39Tc+yuFRa1g3NJXkNMYB55cctIzkJBtAzrkedkYby3nFoUkFz78O/SnVj4CeT1HLJA/vttL/Y
EY69yV5+hUx5WEXflSe8OJjm61cgUxZjt2VhH74p6kXwboMghyifykmhwE762QIoCMmO2WbHUc+s
PzAmK++qsY4gySvtJz/kEVe7YUinW4tm76KEbIkqgOPvXINJlojrtV+rSd05ZUJpM+5GrDe8ta2U
JnUxB8SlpEspnwJ2caemGPO9R0BdaEC2mZR88t8oMZbguODfgEreRVZLqLpIDFfguY85CxZ57UVC
r0JNh3Zt1XvhvDH1WZqMubs7ljFhSeFpPZje9p4krJNac2ULigPHtQLcdCFBbvzUQYFvHNBoSirf
qJ3xxonR3U48vJ6HNI0zeSszjpPG4z1uSDAin6OJ9Xl3noZ0yTjVZWWLcCHNsCfnHOOsqVKeO29G
JsgL+KL3qPRfANicQdSXR2EJxsO3Wjjq+hfQRGiF5npDSyjeI4cdZCeFZvhBb0Ed9tEU8h2+N9pX
OroEX1lvafzqHK6UhrdOidraFg/0gjSyi1jxx9P0Kz1teR15bsa8APDqTTLECeC4QBwMpeOJfHLq
N0czVJ/VZYVbYBpZjMAFB6/HsEA8rXTpFEpm8Qly9xSaBS7WqYIf778ll8OG++aBnKalU3QUMOrl
YqXS0rLU2nC4j1gLSvXsv5m7GWUVp3gvP1MRzbzVSAhvcMS36VhnD6Ahc8Qb23pemiKMnTwxv65o
LMXl7T/jNYw3iJXBvVtQv6qOsAIQ/Xw/G2JYcFCQi6pI7t6VeWZSMYT54XlaM3fdh5W41v5pnXwO
aOG7RjUOfZVCLjc/WhX0Ef3GTmbwOV3eEZRmS5JZA0S1WOn+GG06MOYIVaWWQWN2QSqZMjrxwKQg
Cyo0VKFbs7Sk3vte0y9pTM8fYWO/MQsHXsiwmWgMEmifAsYt/Re2UxNUQ/JThgzYYDyryu7GV03y
cR7H9IhNUQojopQrzvZ+eIsImwLUqdOldyDzoIG0ccbUbx8kYojTaqoAayJxcVcJcVk7aqWE2hXn
s2QcINmIpWbODpVNs7IQzw5utK6V+64kB8vygPVohnjAupNRYcQ+DtrBjw/5an/l/3dUiS+gQzj3
rCTJuucT9sz5IuBoUhSosjZpJOMniXoc8aZ6PPb5LWNBCKKeWvugSsSp5Y4DOGJ0IE2Vu1R76TaW
GzV7aEBo3CgN5byxBxD8DTy0DEA/u26aPJt1/v1cW0VLzbnYGvD4C+Lr0nL1IsfZIs2PoMt3jtz2
dgmeyDNdrSEpMShblTEpXsN1PmUdw8FKiYy+QgThon2B74MAl4zhPT6fSG36WvKm2ekbT3DDnP90
TliMaLvbBY83qz+7pIdXKhsh2wPpMyoI8UikCRkKuE5vAacaYqwucH1dDWT/O8xouIAVNiYeljqj
DdFW5atPegkVHVD8RaAxGV+MaijzPtEQoailwQdBym7fcP3EA/uyMg/NTfwv4EaDWDewTzoKSu+P
XjD69t9lG0vPqH1+/PqFxqClRyBjemymjTm5ugaW/DW2C5tMpMle6rHc7UnF4XlKQ4C2xCPhdGeJ
W/IwWdzV+a/dX8n4jLUSGxZ92wb32ucUbHXtBOl+v3Fqx1O+KsqprUqp8Ts13ZCsjvBtqnohA2vd
VIllBAIf9zGuMuNND+SSbKNfoNx5YtTmFgthiHkZkMYJ1IxG3q/2I+EgkapdOmyqsVf1CIQvFLs0
eX8BWzbzYn/sJBh0uEAn0DlRJbYw3CgW51OzOcrNvCWILXyow8rokJT5LfEryeaarviwRHOn8Tmu
4iPVRh45xF7m7jL74MRXOHCrsKBl2PBN/4q3pnVWLzrckYpE8XxG5xgKi2+Bp6uM25lTw+NQ7p6s
0ZfDTRIdGii9XgF8k4lvWv+Ql8VjMGWDNNLuT5zVoxJiXJHFbBAVVWGHOJuixsNy9ul7HWl1U5Fj
YPNrlTU5poPhvBhrD+I+CW731mmOe6DR8AQuRlayafZZ3J2L+3K9zoI/g6Rc8uKZ5ic1WVoiQyXn
NXBK0BLpu+RpEkBc7jCoJRPDX6IH/Ry0PFE90yXSSRQMYU1rQ132eOKclqlckOX/DQV9O1UAgDbu
v/0gSspKsBJyD5EvwUA34vDiEfGQlP9UqNv37lsTgYuF0yr7iWKf7i6BErlL3+lY4SMBIeAAVgsa
2fPMNNsty99X7/fQ/iEWKkQTqxk0Rlm4J3qWuGghMjqjqEkIeS5wTk3Uz9MA16YICwRen//No/Nu
uYjmtqxIQ5Wq8+EBkIiWvKc0X0nUU0yYOkMPZ7SoljHyj1fAV6QXHjYzExFLc6PoNHQOaZwPYSj+
PBZ0R/Lh62QChx/HeSd9o/MLF/wEMgC1gReKUxFOmMBatW7JlEZKQ/6OeDLeZ8++y4FJdneNZwgk
t4VseLmoDlr6ld76aA793/Wa6Ng2pYk4jFbNG2H8wEYE0ZB1QpVQSl6rQ3VBsiefKFpMl4D8Fbe0
n+8MhSFGvbOqI0qwoe4a0wYxjRLQ83Q+R96sgwexuc+rfsWH8AqMI71sFX62Aye9h790AJk8EvEV
vjhnIL1r2cjxq45cxsrwOOSITrzCS6bDoxjHTx5VNxcqv7aV+oRar7P2jVgVf2Oxsl05sr2cv6NU
s9Cg52gF5raeeNhS5rcuMCwGHWKWf5g69w1Sd328Div5gk42nLhLKW1IpyhKIlrD+7UgB6rC3mlv
SoPlMDn5+4qlnQTJpOYNwZzY+IJllWjDGBBlslux4BGu0pnyq1d8n16sKbJGe3s1JGeE46R+67U+
gNwUEd48F29Pjvsh11ASyTiBJlksF3DQaTNdsoT1cjE6tTrNVzev1XLNCwZNPfQSXEiYJrx7px0R
rOCCk3TOEFG2Dn/g0gAtN7APP/lmso8aoeKOMPRyXt/i1c5Waj9HTWiY2vHlO/CFCS3BLxNBxZ9j
3BKkeH/iWulEN/zKfvyye1PK9LmnOFWuxwBDqBx/We7B3or6MF0ZboOVqF0CFgBM24u57EImdRE6
NTiXi81Z46+/QszPfGHBiJqASr2W8uGdTr2NZ7X6FZPrlI2z8m7mthwA+n5yEX/ljYciaWhloKsw
jWgyGcSy3v69nkczEHRu0jhNnLX2n7xR6V4g57soq+HkEbnidaKTyJ814z2gxziNCACrwdOqDV6R
i4kMgicce2Zoo0R/w5/6dy3lOBLx+zqdXkobJyzV3gH8ITXtA0Uy8lTF2AcyEyVfYvo3206AGqf6
OZRFlZ8c3AoSv8rm7JgeL7XhLb9Qa/glQFLozuI6k7FTtKtDrnNYQGuDQmv59SdHE2wT4EU+taas
1ieKlY8VXn8ICjUFy9i6BsXu2vu11jiV6A07MZ5HvyDlqdM7NvTuszJFyn0WCae4Qdf+5fC7gyqv
UgiFXATGeiJ95hAsIVmJr3sw/z1jFIaqJIXJO+sp5GZBJR2LGQfbhI5ikDRAKv3CJrDMCXXxo9/W
ERGDKLBGpGMVJyyuvoEGRiC4fSE91MKrLZn5N24rvIxIV+ZeaSh/2JslVcpiNgrczgzl0r0noPUx
XeKHdZ8wUOEZ/uW6nR13jvqqY86lfEtydva5qiczcHtla/dMj7NXcWOZHSZkKAiCEyi7FLHzzkdq
pkFXLlazqEdEzGcyMWY0MlWs59uN5+ZVtC2a47fdnJQuisXyfZpjOtPAjCMaGCqV7j9wTLNSd1BP
54OCY9yZeuYkxEpk3lTKYKIOeNVJ6ZF/AFBElaXIir5mQmVMoJCXwRviDy4CRvCUd2AzVNb1x2Ce
/ZfzIsqMba4mLkPruH0BmrOGfxcox9Ph1yqhF/xe4Ihq1gleMUnkwXQgdBZGyArAZYoCvCu+LGH8
2PXsySf2376jqX4Dh8wlBrbPSbJMc6NjbgzC/hERh0okoDUJaqWSFefVebXXi4DbuRN7t/wZnORQ
k6Uxuop2/RkLulrt9MIDaWdfN2j/lZz+lwL0aWomVUR7g5PGcHOKgI6MIsolYBtnYMTSEcjXcY7L
mWKFJyXDOL3FNjcoTYT4eRFBNHcF4vrWGV3ehtXqZcCZBiztIC93KwpabAG7SAbZxUZyPFgAn+88
OsDaLI3zgBo4/dB48Y3rQ54rxNNIfU0a4q528ZrZ4V0FizGzY/v57eFSpGRF0eWMhMoJOE7NTd1q
lwzoVmPEwMlxoay8aSqT7N/+2CSHVK4rfIgvVl3Wjt/MWFhOameTFsVrEuT9cgSu+wZQwQoOEqGk
xJbJjLp+XnYJ5zsmWat9hZ4R2L4Vz5FWfXw1gxWCAq0xHWo8Llca076XV167I9XlM45OzyPWegCX
KtH8Eh2wBcbhTIgTm75Ptjq7ezaqK1I9MhuhKSaHsDjbQ2zCWqBBfeuZSt6U71B9oOAdOLP/lI/v
kwxmMA+ePaTrRfJD9JXau9oFugIWWsFeOMBCR1gTIIWzE1WvmEzc2gJ+hHpHY0MUxz/PUaNFfnVL
FcGR+flOyEym2erp4/a5tluY1gLkEKT3aX1//AyZ4f+J8XdWXkmjRyqbE1FkVmF18kAOmNhcGHiP
4bq0Bis5eQuWt+jZkPU1vyJKvVSJZC431MXLX+zntTIcv1JpUCy5VDS854+DY3nK6x5YWKwAf3Ab
+J7HwapaNTTaSczxZUh1aeoKqRQWh7neu1z0R8E2Mx/9EhfOEahfxUI3jm6dc+qCJ3FM0596t5jm
+lc+Dc7WxRdUcmsUNesH6rnFd92+EP3JUy3M73KnPM7YNySSgk78IjNCuRb8o58Mu6vOsfwLu6TX
/Szj2Dy3cpc2UksuHa7dT5ehCrU36NM9RmxG6FAFGoP2ml1GIs5tM2NXBaEU6wSuPnaAhs+90ApM
/PHRoIsTGUJdKidVIXgczix7X3Gf7vuTXvFXoGOPtxzuUSDzXVy7gMj7+0kGmocK0UjlncpafwKu
CCjm+lqMPi6v+pNIB8/nynqae6vOg+RVTY5j+4p5lup63SpZIB8ZZ+q/goGkEvIvtzDDDfw+z/pj
RYGTZMAVpNKngyrHFpR7o4NbZ7Ju1S0nr1wQQ8b/2M8ipzCzojtKoojkC/USzorFONPnxY9scqAI
pVZcYTRBDQMH8KRIrNAO+ZpvETQ9lHFA5xbFcmVTL/JaHAAUyJwx7Yn0mmSSUmrux9u8QVwp2NcW
uwHiGUZ/HqwPYlGZTxmJm3eQ+aPbqTCL91JWBExXn6tDSUYpDOhntl1DoDPRAHfx67h9CYb9Mqlr
2vMF3yNAb8GAsm5AuEBFi48G0ueB2pqYFWaFl56JZu65VaxXlfUrFKZHFw3g/9TypUxI3i0GupOE
48rKpt7JwbVYKhJvdjtPS9csswlTKSaqoREFo3AMvo2KZO2EVHbP90RW8G9+pcQhfD8rlMu2jOPA
JZR+SZPZsHSGmUzCBgX9cldimxsxhKtlwTpsVYkQp4HKbl7ivK7Ivpl48IYQrNQkj+2S1DF/8qP0
ypLBgNijf0UewJjftqV2gNc2MVQKX5r7Q8etZA/twiKQpxUvB99FVSIyObg93wdksm0k/Pt6kJXM
RC44cKrKTZKQy73z0NxDj3wiZ5Q6UfmKya1ABNHbfeKXEonxhpdhw4IJARm6Md8Td5qSbhqjI+vI
s73b0lUMEdQ16rs81A8Jf92mAf8caDLEZkayA9tGnVmH4Cc7rJ2jCKsc3o4k7Y9MiaOtdJGIxGN0
Vp+tXYLdTK3WKGpodD099DCgmB/oc2+banZ1g/GQ8obXzn+gdPG3nSwn+yQBigiQUzrpYiYkMIMa
exMt3QUppKBUL9hbeooO0ypK7ENcFhPvxmwEjLzw6XVHyJMlXf2jR4O+NV7R1IYggB5xe2NqgJZi
Z8candULgrcsW9PB9Ynhfj4cg8kF2um5Wwxp9Q5/HYGtaEES4FumopZ+gzh7qgCgehhekMRZQRvA
XHjrvnhv7O0AGSUxxahLuC9qfopsuKOczOhDgdV/xOCpcXXrZH8Ov3TxHwd3qmIPVyMwYpk0wMGq
Tjln/rzTx8yUV0aiLNl9+wDDldR2wGCOReTPGwXXkg9nSAEiYEOxXWQym1udX8JgyJj1n/G+Up5e
HBMrEKuLAvsISTsSATWR2g91uN0H7iQYxZDUgrDfpI7ABrNFIrTOm6j160LCp2abisACod7Uyiic
zuDBAvWDkO92UlvmBvSDE2honfIOpSOy0QjI+HDq5mGvBHmxJyY8vJR2i25nTsxdOQJ1BRA+LgWJ
fifVGmPONtoz4zt8IAEp+m3tU18G6r0+QGal5yZ+6sBo25PvNI8AX+8SyiYYWQHbgRSUdjfjNV5E
S3Jv9hV9f19jK7IibFjqF+MXtAMccMhMJVSKnypQsOi0ah1FKnTf+zLJrLyGuzYA6fvMUeD3tNLT
pSHa2IcsQGxJzHaoyHK6gkcAE/IMLlZJ1b37wYnYzOa9Qt/9gV/7a1ElXetrktKNlU3LFkKQRAk5
RFvJgf/G/lvL5ioHWL0SJ8EIQd3fqPjs7KrVVz4izwM0iDBEFqgHKgYTuLdzn9DJoXCTk/MU6Xzn
RtcGZpDB9UwkY4P5yJBAThwHmoHyrGFEseXjmrkFMVFUYpwJz6+bgOmuEXLMx+mrpjM4YDW0RkRK
OOw6kkCBj4QJBf+QqxAq8AzKe+q4rO48RAhqFkw5I4rwVZ4Vp+BiI01iBOa4n7A64ab36JKYolHE
d/9BWmYfHfV0iwAVmd3lwJiYGbeOjVIYDRNaLXV/kd1eof8oI++tnUgK5krykSB1oRUMCW0IpuRy
PAapNMIXaXtr1uKIoROpvK/GR9IYuDQWcz63nL3p9goB8PyFwJx9IUEK3v325kTCfOpOsb7S19dC
MRxDoAley8YdL05B1Bs7Mpjs+u4G/lVOHL6xsjuh+gx+ZVBGbBlYVhLDYCO4bEfW1x1D/9KAU/K2
ZUzhd/h6FW2aiOHiTOOd7XE0m6BrXsb5ifYX1tinMSAE+gNXIGhugw6gns/QlnZMAhkZvD3NOmBn
uURvKVAyr2dIqrZTfnDnBno9G6VmJmqRTHyKf0vBKpWVQtYoj6noYarvJaAihbrJ+u7423x6VY9n
oIa5B04ygjnnAD/0Q/EkU7phW87MbwxGyfYioCWk5PetJiKXcCUgCV5+RpyQbsQ7YggJeh62hpmd
r+3Kyw3/ivcZbCtGbelx4K1XKfBpkB+o/JuQxUXR3TZvp+FBTREki8wcZCnGf4tBYQpJwmAXPpMZ
8cj2LtDk6zXiGs4tzfhI12Md+HAtiRZKc0T5IH44H5S0gZA/5TEkdheG1ZuPKt2MSo5leLBsmHwA
tWzVxC6iROESjuc/lKZGLNAQFDmOlLenV1gWFnlC+jdHb3YxYiyMTkupTtp6CyprzF0493ovA6uM
j989LkiarkspT92P9MKdt8OTfMfoedGUfinMjXlP2bYam7BUm4iwyiI/MHwLTKXUZX370A3AtXSi
+P+GWgD+o8ulh4Nh5Q/U00AUHuVc3PRYbsNKdwwQdIxUCBOKapKex8XkmL6ts8DF5l3+03YvIoUA
xrp/A51yaux5Xqim9ZAc1MgiIhccQ51xLalNQDazpuYe06CjdykLFU/WYGKXkB2MUq1CdhS0zxaI
jUhbQEEmvz422VPqSXsaGr8/60AtD1SRVnVWbGWu1iP05wTJaDNmkBkLNS0ZLgTbttz2g2tGvnSW
7mu7kAs80Ib+8/VrG7eVCi7rafKdrMUu1aTSexle+78DeCyb11PCXlDPVOb4Oj1KEvSNRUG03L0/
DipU2VMIjBXh+J7d1oh5GHRkV2fs7JPm0Ajtx7+uYp1BNH6yXy8NOG1N+dDBQA7jUoexiwfhL0Uk
hjgqhH/BvMZYesNxDYmUABLH8DO3Nz+D+fwN8/q8rdhu1At4P7318OA2UaTXkaR2WMmrjMQN/CiN
PxeOgyoc9mdScSrGXhH76gqUjL1D+lnttceROEl/Mn0v6TiPTTcvVfIaUyjmJK0MyMCRdmN8TQLa
D6/3wrCV5P7upSXveQtzucwZFVzQyYDXRLkEa4ZqD0W/fZSsjEJM0cN9WQPJww+D81EzSWqCgYJg
GHEsIDcnP/owgq9INjPzj/4nLLEANsgdLJCdUYxi4e1y4WAd31Iq6jUPtEdBoj/6KMz0kizgMJ6C
aPN8BbGLG8E0kgheMmPDAso1aCaZITa4m47CuIfUaMHFv4ZVoOw1pF/tv3LWkzdb2hpz80he9sgm
77sDutqIcA5fsDQxMEtdQwPj1hrrzyHXOGPQGo5O0x3K7C1jlaFfKLlUQFx7r7Ep6ohaLjftJ+A/
x3l36rVXwgY2MoPrwKKNQaTZoItozEdUsRGRjQVht6geL6aL5w382NDHx2+/XAx4AFxoRVbtFLyV
XTy1ZXmM0KDbNByOu6rZFgXLtq+O0RLhsfhDIYfb2189+TDqIaLQDLHxps+wu0SNetivdHYyM6gw
f+xtwPD26Zh0tQiLZ5R9VuBmH46841aldv1dPN+Bm1eDwiTS03eXGCSWhuWotSThhpLxcqTO1kN9
CvFUGYa5X/YEym8x8xo5M2T8D83Pi5hRSKL0U0Z0APpo0K7OKSKgUuTRonImdzxKH99D1gOqs0Eq
5BOlnHjIovekWucMLMy4dZc8lzevx+7j7bQ470G0nNMq6l7YOVfzOmhJWz5Goh0tBgajTa0TweUk
Rw6lmuCXk/7SOwhyzSV685FIBKa6ORZvMN6dbZKhKcCkvhyXdUEi80PVXMXpo0mihY7GFYLgQXPV
MKriMAoIPAJo/EVKRzRuE0O3ggh58OVzzMi+0lKqBriVY8xOS8TZwJPjrEVWr/IMa/6SM5IGttQz
fTh45idplEGbUC6X6I938Kx6fxMruW4EVBNzWy4EmFmio2vI/CV27x67CqfeHIqrT9qxpnwBLAjb
tmfUQ89M1bqNx+ocDtTdIIrTRfKHNpZGk7RkUdP/9lOc3eUjXpyPLNPACVM3xwlsdPquoY1ise4n
a+y5hoCpTHNpTFgpNIEdmEtBtMeAqxjjWBYNOOCYJ0ghIIxrGoGw/xLeDCifXZ/o474Dkkdbv0ht
/IP2Kx0Vh/jqXQK5tyLZifblqUlRi5fjDmAd9M3u5wzlCeHEKEKkqXlihmX5keijtEQ73aCP4pkQ
6xwPcJjg7JrEGMpvASHUvEmwrSPYhI+LgXoOGxjPgsSMCEYlkDj5kC/awAEhXL4L9/vyPB4rDI68
rgPj9kqkZZcFuMTCkxdnLqvuvD33AYbf+tpE8Thk9hJe+PISncJUW0AJE+vXGsFUTnsVf9+7zHmp
Skdp71c0TfC25b/ekIaIQ+nVCleM8r86JzBfcKCKyvrZllbyUdBEbfSxvyK7WArCkf60zGa7BonZ
rO5uSk8xw0slD7WeIRqux1tIC8aYCM+evHnIB3Taf2+6qsINfPuKD3dYybaBns+Ydy+WTGP1fpuN
sAbGlAxtokS3DDy/cX5AaVqcLGZqkTGZviKsB3XIdWU6956WAilipS1cwTUiO5DACbk2SJDgsB32
KksM0SWa8BzyO4rWiviCf34CgDuo4F246Tvl4KKSrwFROuiKLB4YGlJeAkfJ75fL+Wv1Ex/R5vDg
TQv07y0h+TvaibuDkh9+M3smG2h5bFO6yuYcFhRba675GS3/dF31gWQgv7MLLz5yU6tvHSAbcnH/
1F+UYcw42MXnpa9mU6yWCY8CfxiFrcrcMrZlp9dWXUbV4q3AFyt3GpohmyvurGlnQo+FANj6v00S
xw2iY0fe4vcOBzQj2cmHckCmzecY3U6LLKJHmUZS+qC7yYTYrejZXChHrTfttOLH94hAkyVawuu4
gA2oIqbLX3aDM8NLkI+MPc8hggFHcZe66Iobo3OfC0stG4KrfCpHv0fu2F8nxmnyARJob/0DLYGf
wRIH0icyJAtqsulS0bFWL34U908IcRoyFU6BmL2dcXjqfIuUn4urPkhWoubDR6XKOy0tikAjhCmg
rVu6hjlOWz6VW1QyNRsob6CCGRAYe4uWf0YotFz71hIf7c1UlaM0Pd40s3S9VcJPQ3Sd6wUY8a7d
KJkuOEvRnRrEeYW+F8xIWzuEF0OT3ZvusrIA/FuxU0ofMxb5aLZ3RseGh9HBvoXI9pnSeV6QVlAW
5Bd1ZSc/vZWFHk6ckwZ5W3EFgOlY5ctzJ+OYA7D4NXgkTJcgytBmogGI4GCV/vesF6uJ2OXv/u9k
YQTLg/GPnnLlwWjeaZiQwN3fObwB3eeUGJ0pFMu7P/Y2/u2c0BeGARE8M+zKpXLqsfG6ILh1jku7
kUF+s7Zkg9dErTNq1lurOz+1T8WHxrtoiH+hr2hOYufZQmfAGy0pnypX15gJK/2oyonnXl8Aih5P
OqkjUD0K/33uq8mUVtwsNUI3vrC4jHoIB3RZpgjKtoXztetSbRH2+YSCKNfDPsQWrtLFxPo7kZTZ
OgXmmg5NFix8eQiFg+FMhIiQIpVzAsG9TADUpmVa5CCuB2ZkVHYQ8LTdMmZCG48SMLzTJ+iN/TO6
aHtYPVM1aCVzC9y31edxOi5NPK4lb3XyzsAgIKgiQujmrYmGjCmFJPkShcCbRF7eUPKQc3O26gVK
tacbP05YNcJBgDSg/XBCzlbclF2JJJW8JwDk+5ReKipG9AthrBdF+/53r8RPPrNq39McEfmSaGLJ
xUtN8Yi6/6yJk/DWCJKvab4L5WV81sIX0brN+OsS7t2JbChttqKtBKFRRfIEf77tRu+Raxge7vAv
ZifSdg1XMGNlcgKtO27U85OlhWqDWinFlG+0uMh51caydSSiVAyL5Y8wsdrdUBvJGJtp2++Zj5Sh
c9zf15LWNpWNLd7tMRO3FgBW8RRP/cEdqB5A22/JaKa/8WO593HeTisTCNWS42CCXv4M2tgvgNyd
+hnHysxH/B0BDaNajLdiEfhxZRf1hMELZdAbH4OIGuado2ToHTAUQIB1PAL3T/5GhNtCq848QZTk
kbD1vMhIcbWt25iuWRzHJ1ogNIj9YKs6/q+NqKxZmZ09oBX8rXBWuHegBD5ELYtYhOxoP3xebojW
I+gHLTX37RMi8rClZ5iyXFjR7AFkLOHhAa4F2kc0+j0WoHbU8emdKZezm8HwQAHkglWa40hdyq0W
wsemm3xthXt2ZyTc38vskj33QfWfy1Wz3AjxZnZ+2grQERnsF0MBA87W9W5kXxUrTwrNhL6xGNKV
DJj/WHf4Mx0HjSRuFxDVsAK46zvR9gtBOyKURcjaI32Fk+X67YHgKttKiz89OiuoSGtrtq0H3nxg
zmsT2YjXL1QppMVuPmtaCAIlfKT5kayZqY0qZJVlSyFpNYqNojBOUuk9HiGyHV7N6T3KmwH11t4/
3nmyQpK+9vyd3iABBqH2+xA+NDGtPQVpVzTmKwH9CJRd+ts568gMx/FhHI+v3fV//uWRcyUdqaBz
yK/HxH9tuLc7dO+u0RIaAw+kvLu7apjaLhv055mbCmT2SmO+5rAwbolgT5FCgRstTx4uI7lh2B5K
Icty15Ws5JALetqolUlxX34cUVMVVMQFU66pJ+E8Qru2FOIfHJkTVDbaiGJZ4by3AFKaY6lfxJS1
7GHBSP1AojrbbX5l5KazPdmA9kwbsszryoIx1pMcRojoBNgatzGVBEVOPmFMSvoIkAx/7AuP/7FX
kAFXKzb74tQxlBy78ZIc5utTmC+shKVWRmUJFvcvJSC0hKp4Pp7Q8a/jz1AX6OmgdJPqRW8/4Ocp
K1vYbpvn4LAIno1j9f8Eqv4EycPZa/rtW/4Rik/yMkzS1yqAzPc0PK5CZlh9o0r3rP3DLEDkGxae
oBaN4LTy+QWb3beBwQYVb/seVvWq/29Temdkni5mDg/C/ImKiYaKzzBWdHeonFao+0aLfw6XllSx
dWANuyCEjW7B2q5lNeA8NbRf4xJ5ztxmM2mqu3gMw0j8gONL96BtDd5tehFtgbf3EDZ3S6XM/ooR
dQFNX3/hVRwl0wptNb0zn1CWcSV3QUQpVaKJAlwBcZNjGVmH2XA61Ath5r8LZJuwIJxm6Wh0rZtG
0pNgdKHTwgpyNPXEOriqAuKuj6e14JFqER9tWar6mzqZprKSbfZJgk2oheOqP8SWgb7lAjEWMJMe
oAnzoa5N6Cf8MAou96IcuTlXd+B5bVCUYfVswFDv8erwz3/96r1dRFXCaM/iYG4n+9caj5+P/3I3
gg1JZUt2f+4ktJmGzGufwyAndQf9CYhmQSKSBaPn7Zlnr2iERqihtfqylJQy1bMalU9FcFQJw3sq
J6zNnr1zhgB4FwYvaEJKv7/ZRvbsqJUiGN6qd7pS23q3GddDDKwSFgNG607OqxGlHs51FH3Ms84+
LRL6xBtQDYry612rBYm1i0yhgq7LvbYLrgXOlZI4Nn1ckXws7RadtRtJXXa3G6MpgZuRPM2+Au4V
bGKSXLhGuWC/6JAjMnufGD+kMXWV1XBJJLyngX8n69XHSM7yUrBKlWmFCqd51r+BjC402FF3GYbe
IzdL8ZGY79gyf2s0qeJ9LZcWCUAgHhwm/wq8viJYPeCrnce5TbXRA9IawNlMj/nxVP8tVMvP+5kd
1oAq69l/CBOaaeNFXjrZFU1ruo9OK8QfYxADZs2+1x4dGvsFEFbygtFDF3K7ki1c6Pa1oH0/56Ie
Upelx1xxOr8DqEdhv+DVCY/AfFalFt4spKCmF/KAkOGCmTpDELbNJDyy6UQEOCs9T52uUpyaPHOw
NiUoVCCkwtX7TS0UD20gwBz7KFzPaVgLozlLrvxTa0rgRIt2Dngb8GyHekqEmSPRYdd5niTQZ8ZM
USLWEVe9BUm4r6CKNr2wYt/22OGr2zAu28LAz8q+nK35cTBwmkcF2t1L+gzQRS4QOsRESmuRg/XZ
ESYrA4S6QZujK0lac5WKwd9718Dd5E6L7cEVJKirc3WJgRCFaDnNz4pM3Wlo0skEBpftorV0st08
zOskE60bPe0wYWUQqu8Iw+yqfO/8ylDJaloIu5KYXgAftF8LpiIcPftCGaPEYMOzV7BIJQJHIwjx
7oVlIIuWuslig8Gw4IJ8lb049etjIiI6F5xxmva4j9quy3HIZNkTJtYGztcq01ohgT9mSCraltFv
Eg+86ouRXKBP806F0QLzmZHq4BFzdlpFUzIxCdFZN80sAkoXXqn8d06yKUNljLpVDo5S3ta84uj2
rcbGVLzjw8Ww2x/oJ4tfavhIRlnqDN5G3/sNKMOhwZWaQq4CzjxJQJ8c0x4kEkf6u4ZTThSYPZ3i
1L1MPOwzfzzoqJ5w+pd8IDkNuT07gQG3FejtmSCQ4Se0/BB99lsf2WAwHNjQ4YXAg8lHbJ1EiAam
z17Gp8eK71fJczKbnclX7YlZIyscBDM/L5LIsfTHlmWM4JqwwHsTx7yqMGhEgAFWYI9TyT0AljpO
PZHzg0QEJisHLhsFkU9byg1ve+LndZLVrAfEK6gG1hpex+8MrSf/KPo1aCHQDCnxrIIHEDanuVIK
bX2KbA4xLexJGo++pszzfvI9CVrsuSUeUMTfrUEEqXukq8Fc1Jd8aJJ5/d62tVdlnVckxupfx2pS
G12Dz/NdDi72LDtNt2fRZzYUApWlw2iqYpAKgT9V77GMftPTqk3G3Apoe6MRQUozUhmCXCC65BGN
iYNfTV8wT4BVOTKqHUJbpq4fyEd/f21M7bmTwsryg3JRC5K1ji+LUPngFPgJ6IQBWdnGH3dtQUAQ
N81Z7Yfq/KMZQEHYQPio9U+feZvwO2koVBu6dkkN0p0CsiiRgCGDlGUMeHGMOUBAzectO4rpHDIq
4tEeDtMTj8EwPinWeb2/MZ0KWf7cgHKCBi7ycV7odtbSVrtR1W1QP6fFh1VKWdMNQ69GLgVW/Wzl
wleMGo7UX6npVRZ20CuTxIVsJ5t7dwMplFbI07KEJH96zM0aNpyeMvyHs+aJY/AdRe/Rs9o/PLhd
TSYkx00iRMOZd0sfPt8BtKUbJYq2mYAlitb6T4t9jxTjmsd1j5tJX3Kns57jioRmUPtaSfDbTiPb
ubwktwD1xupTF7f2K51/EQ1q4y29LiwasTBqaWgGrFocCRO6D5qhZ657pQ6voFNH5xa+DIgobF8R
2S3tDrQm1szny5rtiHt+DX0OecqJmPu9X1/CltQixIH3ZTcI708KZlw5IWnxN0gKkH+nlCdjIEfd
N3lfJzLaXPHJJQB3Jt6IR/FIBgkosR+8EXvimOOMNcD9klcTotoD4fYwnBe63WEiGoGObpw4Wqx7
TAkfACEbafj9Ds9eoWrDmAOlfoi07QbEr0zMB8GjsZbwWck4y+5lqtO419pt+6FNMCHT52pjrtj3
I5brEZMi+GWHEkF9YTikGg47Z6roZIEJSgLWESfUaZn3sLgRdFOGrswoDB7fuuIivKJF7glVG6Zq
xTfKAZdnSAvj//mJVzHk2StgISMwQK92uts1EjyKL/PPk5Y/91Iam1XM7zwvGAuAALQ4BfDDjA4b
oY7o3z1Z8tprdLRqkZ3k5jjrG8FvMF1cJb71oSAKFfFZxDLlh2LQGfzx5Mjjqp1qjnouiiqIs5C4
Z4PkeRK9zB3QrIhEI9LOZqnu9ktVftR3FcvYux5Vjys/qgyBs5GDqi1vL/vqeClxVAbWk86FNbfo
H/qwgQYAZE+vNB0jTiLFkSoOmgcAPe7SNJjVIy4tJrxpLC0E9wAdvv6CtoRWVf4/Oh7X5YWZch1R
SpJWY16ga3mnB+VdquKI+LsxrOQHTqh4EczAa1iDyQWs57WhheXvmaTo59gV4nHqBOzoZmBkd3tK
g6fpTvXHV2ER1IiY5HjOen1oWdoxDzmYh8FM6Qz29kTmEM86rjkkFfjDmH+dSBRjQHi9/dLnvwSR
8mo9P9hwIyIUumMlYwUdQ22Pg7lCT5ZBSZT2pWJNPlf2HuSw8SjXCOdPIk5oSdvjB9UhSUNENXI7
MrZon6+1jPXahZQwJssmfgTL2cnmXUZ60lZcAYbRBXxRsrNTgI9uF4kd7Kj7WhOM+8EV93a+wHgT
EnHIsUWnklrW16QJcLNCG5GzD320R6bKJJX+/UJ0GDV8Phk6JY+YfclMuqIWpxa0gGWGaWQNlY+m
AxlZjlk6QKbLuJC1JMoT9EAuTDwJwCiqlLd6sRHcTJFw0NoIOlRllH6IzPg2HdumFjNChsuCpHyy
sp+tS6Dvyux0+Tr4xkp9N0yEFjBPpLNpCjbG1W8qfKnjQ+X51m+xs5C+bZ5ls5y8iHauqPWqX4gr
LF1bO+FTt93RmC9GcKURE4Ftpj1Rc/eUwO4sH6G+H2oYykjfSGu8rAmSrGIV5GV6tp48rn2NmGgl
57UQ5rLvi6Ec53BYZUJ0+7rjuuPpF/Mz+VKQdos0+UJxhkj0mlkCaGSH5Ez3SgT30a42bINphRMC
w/bbWXP8YoNCDNOtAugn4Cvokl+g+f/ya9Y923NL5eEcaAWiUBMXaXcKJ1pmStbxvpGudWL5NHFu
UC6IQX3bZT7VNJX9XxIe6oocjfKxeL3UgfS14gNinWAE8jYY9wCu9+9Hz80ZYltKjILE9Y8dLWYo
L1lHuc8kQ1sN+yBEgyUdYkEaSct24ZZvXi9Cc3B4tNqbgCBgbEP0UsNiJ3ZcxiOmWXqOW8s4RXPV
tCjXykdSHRVR7XW28cKoTB7KTS1BHGAlCkz4aLdWIArqz8gAjLLM0JbDLflGHOY19Oot25q/mNwk
m9zJhVGqJ3/b+1KdP1BWYtizVUF+mm4h1vY+fny+76valpo9woduJ894XCN12+Gfh9+un3RMGlJE
jWARfmUWarEZ0ZvN59vFJQ4V/j2YpnqM8mAVrLbnEbOFYLlIN1tu61Nh/VaDibyjsg6s7H4hR/q5
82VR/Jiv3aNNYxoLKP5KjPe+T4kZ6Xjq19OLwAEgJ2o7HRhR6OVpi3uGaJ9ijpAQYH8SjYzUueHl
tLkZVPHb+AGXyDm1aRhhTpCqvkAdrqveb7+HA2UR2soSnk7kUNZw3JOFdzx/E7YzjRQfj6e1NNZH
53pY+wpxhzqzBTRirg96gPYpztX31c3e2KpNuPVPqrZwC8jcSop70TRlGhAeITjlTQ203CVrvF1X
JJvpmoDiT/3AETaZI5cSfn3PIZMLeyp7IeHA+aaY40WjwYEcbvp4OVjbxuQclbRb+XaJabairNdy
Z/tJFtVK8LdpiTWBgQwMsyy2qyaT85CpdnEDhl9jKOsP0i+axGSIN9kpePhCTHKr6gGUUF8p3i9C
qGzUDv7hf9B34Y/OhGEhCKVglC4pq+E6YbS6cn2jHfxQRIKqmZ0FBE5L3fGvS3wrpQgBxEm3GcuD
RNE1KzpWumdFm8tSNpyHwHRwVzpObr1FATaURSStxYLYxLYsqBxn2BQtP/kncCjc6LwobuAF2e1v
0WC5RYhqumTPVYpGuBA0qaXcT7rA9hUg1MHpO49il/zYUSKE9rvTi5LZroZ93nH9cG1NPVavc4Vu
8m4PQZIoBQpTc/XKc94XZUsQlAlnD3Gvq9fCfbl0oPeLumN9dNWu8in3zfZ7tKv+euMiFp6nL8Ub
hkpHm8x/eCNY2A87uqyFguuRKV8m5VhZxsVlKs2vjScaooLSfYtJhcXJsoKlFZfmXaC02q9tXKhL
bJikhtlvIp7O8RhiJgBrntZa+eQGJn67tIdWXKmyyKuFucYYU3WcDzHK12/LThYMX2CfqXUiDqi9
8fSTacmExmtFBuFor20Etcqm1WvJ8vc1joNdE5IfGxIv20W7y3HJJsHgBwIHoAP1DcJaMW/VUl7n
lkV7cWfJydPqKTubPvyvX6FvnO5oLEeaSWnZ9SV9vpfWFyOJOEuzvly80FHt4VgRTxl7vW9W0lK6
IuupBhL1Fb8BRXhH+4CYbTPd4aJPypA7HrbaN9U2PeiHqZFLbFV8CvOkG6qKU1Tv+UiWal0PQ8j2
FVqJdMxlluN93GZH3VMgtTFE696etGFengr6vwONWROr5fsTdU1sro/EpMPkcGzv6lW7xRZEYnFJ
K7WqLRKGr6FRYNZWp6hSTr5jc/RkgTTy1B2thX0q43txt4cpcfpDneUHOW7Ni6aD+maLSjhviEMA
L1mImwfyUNWy30qXqmCQanzGGi4VP9kbPvxM2nNEEtAOrRdLZk0aZUVWnpbIKSylX+KRzXZBq9V+
wfS8pQFYmXaJuoMgqbp7pWA6WkJGutG06N/QQ5514on5A4fnlYU6yvI58+cj2PozJ9mCSP5SHIho
dab6zldDSZpFzbeFeR2W4fvryOPQweNxoowfB0U0RaxMcVF87k7c5NkL9xyjvgZx73gMzO03mdwO
tiJB0judus7YtAsgoAYIQkXQeUebEf/GlTOxdEoJO9K1/ApvCPodprBgiPgH6/W5gLFkGqiHcE77
2VzKf6f098tUido2+2bvGnkamvUxEoBYSDPiySS8Cab56vSJqeTKjXb5xWMAYYAWs2NxRS3Q/sgs
Ti3Yq8SztpiFcO3opgbluCoB/oCfM0ESSCFGz1YubK3ag4AhKrvagn2VyEHolMozUZvzdq6iQX/7
gFJVnpxISNR+xb+9YGslGUVAIl6DQ0sAtoGsuQnZL/23BkXifWWRqc1mXinNC2fsWnl0iyNl5+Oh
J+aCIFDLxmdv5X30hnABEAFsO0lj5E1r47dvpX9LYLa78GWVLdB5bLnVf+lBx7G6PTZ3ISKwoyL0
xfjSd4PIe4I/NaFESkMg5aJX3iZq+dL4/K00Sb7P97yOxcqDeE25aywmLv3JJrwzCsxJhYCAM4Jv
9FiC7AZpDuITPBxgO6CxYUw+G/EKgQf6ThFy3T0SwwTBVE6gfMPKk4CTqMUVPXro9dgGFfcpmaln
LRwODl7Q6NOU66mTDyId8DlkjlpjpJPYkGjI4nYwbgRNTamWtFYIGyacASMNmzgBQ2NLntwxCPMK
s9WUbOWV/noPB3wtrmGLHVfMg+8CNWJMaU9eCSnzh8f80xwUk9CFdmGmo4UFn1e7uhSeGV0xdJbX
HGgnYRoeXatCP1G5wQncwTlihBsUEfecfizb6h4KL/GtJupqoIBImq27WD8yJonI4V3s6WJX0nBi
hIDcnh71QzoHId00A19qNJsn8Ez9XRd9Q9GImss3iILVhNwuxS+rB87xerIz5nixQUwVvCh0DZp2
157AnVCs1DvLNLvmVs3Cd2u4GqgsecIn8qkGIxkAHW914CRMbDmubXsuvM+2xX9lXpSmD9K+vPmz
0wVK3UaL7xJwujic/3YAC54Cr7g6bZgvbaYiUrUQt75WoOwN0tjXn3fnMJLTGYuR/cdppUVta54I
Ju54sLPcKXJM4M2lYn3Rq9nY68zAE8xJGpLsGwaFpJdhmnZLa8cUyG9QKn2/WtxfU6XJFzp0X40E
i+HCp2dwA3jb8nNM2t/1zCmVvXriOn7Xd8qdIpy2UtG0b0mAjs4V/ZN/VUqpVEwdoRpdDkTeax6c
C7aX8oIIliaqBIrq/cUGrcsVfZH9CpwyqEvwBVc42v14uz8Kf/P7o32AxOUzXLyx8EqFnnn23ED1
aUMXWjYBIS4Cp8rJIqbF+sQCVX8BlCv2qKFtUNNwo7KaU5qsFY378PwCmmY8i80+ZjDVy50PPWCS
NzGR5KpaD4RA09jN9Xd9GxfB+gDi5WsRLsEVN+rD03gwLy61Fhtpct3UXpXNOzIZcBBQfQbC9jZu
cZEG8quxg8VcCTdA+lsZORCb9/goCVE3bPz5ljrjbaf4xB4gBT83mV/leR65vJi+4qyBW2DKSybP
Ro7nRtlz8mE7npD2pBdJN6U/WHdvvHg0x1ZItgdXzwyuzZsGPE06fXf+MDC/Mw+2TUU25doUwlrK
n8UoJZm9+fOsw4sZNdgI29ZP7EmZKqeYQc+arTwaoZfGgTkYKcL6Zjzjwj54A3FsSzcIRmEtCk5k
wE2jm0LSg9FRJPeQac1FxNSel/VFn5ZDkIryPvoDEvgFPa0xuaUjVxoDexwkW4xL8Z9BmyIxctbm
IC1NuUpSiVsx7ziOqGyLu2NSfQulAiOb2/5Voe1nTO50DV0at8AeEWp+LmDzz4fdmEu5BbnGcTFR
c/qt7ptUkreh1HEblalCrJN2+WYcqz7TuUysdf4PorEd0bkClT1QG6kiYQ/RYmnKCwYZLrjp/cIm
e2zDDo3CIVkc81FPOtSXHsgXgD6m9MY53U3NHPmFiONNV/MwIRnmNw9bv90w95IcsH3XqMscs5r1
kAxEDVxe/ldA1F2nlBIRFEwsZnt5slv7xW+LLA4FyqDuLPgaZJZlK8iWgcuTZvBx5RBQPDj2BkRr
tvHmXstY2+v8GCqsdCTVjHd37+GywJdgf/PQ4TJkYlwpY6gN1JJiVB8rop+qwtautYpNdHObVUbH
eaiBeOlAJ9KQn7MjQg1n8zyBu93gnJuqo9qMKHeT4y11lmv2kkQbmYFm9S78DFBRe9Ix3n7pRn2i
o8WbL+nJRO7g4lQK4YcEHF+E9aeEi/e8dSQVo4i0t3suuHRNwIw5H50sEL9JQCBSzmzLF+Ue7DrP
6WRZd2ItL8YtsmdSjMjDvBF7RKy0+yf1Q1H1WdJNxKHElrVxV0Y5D9DSf1PgFCKrcRk74BU42Cr+
FpLvzH86ZTGtWV73L7Umw+tvB84o1/zSmwqr17ewldpI8jVvbvSAHwCUMQeAi2PWv1Hl5pM+6fco
mnsuP3mDQc1nUxmNV6IScMJr9k6BewOxlCUhYoC0S4DTtVe6QyVJhOB1jyvmfq8Z9Kqsjf9OIv3V
VHoHFOtOJO2KKL3TKPFdAy40IV+C6aUV8Ygk3mnwNElxJ1QBITVqmUQX9uOe31pfpBmxt61mEr4F
ThiBYsC25Qfh6Itz7GKvbumtG32e4dnsfOwWC/sDHd7W5Og32MCQmSJghDIuGvLm1o7DjtmIjSq4
sk3EXZlbhU4uXKoG8gSkJ4lueRc3O2yh2Fx6a5vdv9SB91ZsfQGqWz7yTPPA+bnQ55R5mvrapbK9
Ic3/ffQdTMm1iSmfDuvoB82lpC9htuEqTCwxufmkSUGWolHa/XzvLkoekBdFS58ANaMatSswMtF7
66yZz4hunhzm76vGD9uLbNT+5KuVF7oGhZTGN1bk1LyIsCNIFV+QMT0iOt3suJvnzwyUMYDYtWy5
myynrXftINJhxOXgENC+4p6midW6fmiKKx9si7TNfenY2honn0pFkZtl+CVuLXBFcXzmRWvbcjIY
QiWdDjfZqxpYX3DB7RO5YOwlNYN9mwt1DmzrSrAczPBX17kzzPO48ewTxBsZnRg2u8ADMB8FrgYz
gE2Pv2WLj+1TBE9kqCirlAuZJeTzNjvKF9bRN/Yt1iX7Mbf4bknWtOAyLkAewjAU+toPGye99NEu
y3QX+BwP8mqIdDEJCCoPY2sXuBdcdSWoKuwS+jEP++ZD37AK7MYeRuhMUQr79RIYh2PbAunig6Hb
l55psKpXNTM8jnhC9nGHj9B6qeOF1j8zDOX7Wt7QlUNEg34Tf9uvMUp6G9UVJPOuRc3384sDupsR
OD8/kzboex2kA3Gk7gl4zVtL0XoHkFv2dlICAUiKQdV4KRMaESDfUoUqBjf1eQqRVTipU2Qp8iW5
gOImncAIsgleBXcWFAidUhF70A7sqJ/bhyv2tdfEjLk9hZltSfTNNUNDOEdYyMEemkJ/LF4WV1lM
W4F2MSYPYDlxItbdV1MGrZpugWS2HBHGaGBQ2n96QPU6BWF6J9OAHnDA63v+JyPpjNQbH/0R8pME
7/hY4TuxjzG0mE/kW3wxvsMzI0ZtAEJQS649qMjqooWeVva9ksy568alDXhOK2HAqDeQAQwtqMQs
EJaZQ5P6t+qofyOvSE/FzoNH42d20HGpr6jZLra0PndRYkeuGLb4ANXO1uSN+V1TbJdUvOfuXVY9
BuCNxMketCPUUlnC61bgXILjD+MHM0VgJricCmnempSnIjOSU/CWhuaxu+x+QkKTiC3kJy9BNv/k
lcLVTnjtt40v5bPM8PxmBvlWISJj4gi49kLvS6Lfqp1GdkAQUa6NmfiVndO/BfOOzXUyEdaW67r5
PaLC5EZDj2U17HmZEOmDPt1/6905I/BvGWC8puVNiokVQ/llWBnnvHZE6fVcFXn4xR7rdU90dxjl
HlQ7FgzyZ3R2OZdLvs4ThhXHnamrnloyOLE39ibuNWFB17MBRlS2O0bwXqQZ6cEEuCVsmGqG9qkf
38cZiLThCD2ZMBhUU1kAg8/NUxkX99i2Ze787JHL5yoZwfmuUWjDXtm6/sJHc3BO25NUimacvP+V
DFWIewdTeIIQAtfSri8nnxswLy2C02Ugj9yjxaVgtTwtAfEFvUKJvf58fZxVQvGhSCyDmd3Db8kl
Q+SE29/JlwyQT4DMK1jhFycFYsVosBjcINTvv4pfNZh5OOV7GFU+wY3fIIXfLJyG/lnebOZV3gaB
KCMne1F+NUok21E7aCXBoGm9hhTMRgSDyjBIOS7JjwYgOtoOssxRDHMxQO6yHahCcbCmp3K5F7No
FKbcBkG2i6RCpz2feV/FGJOMHy9HLx3IOn+0EQ3Yuc+woa7vRkfLOq9Y/SSZelYUGk4G7kRHsoeK
OyKFhYdV9sKy2e9RRZIfoq0M1URAVIU4Qoica6ex9MMVIr80W3o3MjiHagk8bgcK26l7VIrYu1uD
0w9ej2wPfgl9JMKbXpi9qdRMuenb0OQUx+xsEn3r5eGgFFDSspJG0nODohPkRbjoIXT2r5PSSIUc
e20Z/f73YaPVp23dwZiahdUUpJkNEmVohXLbAJQPaXQIe9ckDnytSM0xRKLcQLaGz9QmtENcFNy5
phP41HwzfWB7sM0qxcrHHX6TRLIP8AKbGexwEMzTUXhVKkAXVi3v6uECdQG0eZX5KNWaD+3GIliL
KC/sPy1PSkuS9X9vRyz2QNTlMHjvCueA9/VCMfWMxa0m4xxvf6De6TzhMBaC1QdoMcUUXs5Pn2I7
P0k7Engd//efWFCT1IhXFKoi1sVhwkEJ1WJSGMw1hhwrvcozRDZoUiS7alprEQcibo1PDhYc+eai
E4ve6vwpITxFurOKlusMuC5qAK0Oy1PWnd+njAAI/Ung5upK1RmrbISjvO+Ob6PQg6NmYz0gzua5
wHmKL1j4DRJ4bM+0FBtJaUuz2mX9H9C1g6OGTj7tfCqose0f1Np81z9a6cDszfkLrUfX0nX1Eb8M
3uBpw93iNeujsIArnzTnWlimS2zAbQWf1FSbjvekGV/ToS1fMfijGmpKIT3tsjsVu87rq/i4sQDP
Bi/t4fOO9q9qQ3uo2E72uJ/RLTdHjHPHvKRr/2IPhJ4NHACHkgDbRFhK/WxzDUN8jpVm2+0zIDU8
y9JbkLNQMMMrFdi91KxdUPWdR6D47uut24km8c6cWDOFEmk9aky2VwUDo6h+8sFg5WUXplVTEhou
tvuN8hYumKUKP0MgCKFwvaYjWNwzpuycb8oEaUjmY2JexfsgYUB4KWd1uCp32tIPSRyxSe+f592t
9YDU/7w3ALg7yQ+AaQ/Rj/T4vEiASB31TTCx0P81T5QTnd8UOY2nkSDoxTO7pNh5Y0Ole4qIrGUj
kbhCjNOEH8IBAiqjqyjsHosAeJBwt4N6rk/caMO57jkp1kZ4q6BYP+swj1g1HcxbfG2/r9/0/b0t
TcyyySRTHWKXAzm8J6ImUyUYuswTTdJHvgT+QwtddeNREJU3eVm+YYvsJ+pka4XVuoCk+BgO2alQ
2ojvaYDW/FYGuzd2+ijXmp/abssZraOLwSu+wkhgKvAEnYBeRyLeCa7Cu3uBpw4+aNGeWtmPNT10
eYBIDICWvo13+gbYeEzOtlm7ZZmSUbiGRfO+mCE8GnZ1DMKscxymc+DH8sWMZpA+MY/DslJmQZqj
5CAeCZFwDXqZflSXtEKV1Nl1BB+01Ycl/BIcVaU5zfCtnyKegfP+fJPMdUUIgXOQUERPeZwRd1ZN
jJlIQVU9tg/D22J+HG2Bi/3JjOfDE6+iJ4iDjMltKr5v5n94Eu8fFVFgennK0Nqfe1bCWg8PYuzw
sy9DLS3PnfEZ+yXzkX0oP5Yp8Gq1IDpjqeohadBpTDPXN8MjTxc+SKo4f2cjcwswDFVsk9AAHKz3
VZqPZVsE9bjWeO0z68n3nBL59xrmyzbqdQFPpPbN4CjzuPFnFPRREuxsoSSb1u4GJwR71R7C88f3
rDrR5r+19CMEU7Jo53EBvH6UKw+r8P272o/wTYqqFhZMrH1tPr1jBA/kM+BcG8Sszpxdr/7CnKRy
8O6d/fFFYfNrLXZJZc559x7HjAyoyHEuP+YysyIlZXSif/NDrOEF+xj6bGJ6A8yrX8Y36mg2TDdE
PQqgWR2xi11vjlkja/nPekbe833kS7kuchagwlc3mAVFvZlclOVYy6q9Gn+vt1snUYQCN5D/Ym45
rwuL9vjWBaSG3BYSE1FTP10UdEXFUvTQIQaceCyrtSk60tKPbAeBeI2psf0v2Dr7tWGbdcaY3LG8
yZIlVF0XdRcUnGuYN+V9ihUcpvShYdn4iieupTzZUonjE4oBTUlU+h3dJUr1SFYvSAWJ6BhD7I79
ER6bju7COy/J/eYPY6hbTbWtu4XC6s0bziU/4kIxn9Ex88dXipHFUbD799pYP4WZtyiUc50gQKH+
gia/XGvQ/sVv/IAyafwBCaNdwqN2Lf/E+4jsflX47yZFDYJRfe9/wBYjt5SD920e2Rzh8/rGbR0u
qkFN5xlkGOFOrpWVj3zPnLF1ut3EYzba6G51rl0DOQVuo8sLXHvBIxbmm60PTJ0J/q65mtScmkET
T/13e45IztCqkxa1Tb2NcjgNMs1OM7X7DIErl1Q/6IubyoTPZ0TWXn8dVWDUuo70XOLJ6M0Cl4NX
J9qx3CNxBsJ/Yg/QiAQTxW9JaU0pQWjMNysp2c2UwbWkD1UBQRt1nh8YDrpt7z4IKkkH2fcoLDfm
1tZU/qY0o4+2D85l/nETENlgDuqFNO3QY4S2MElOHKVhpUdFoaZmRNTdc6EZ2OKQpCm4KojvqaZC
scECJQ6UUQsu58HqJFZP8g4D4Z7V1FlBi3ArRiZ80dxnag+1PP8JkFViQsDSDtnRn21ChbjLF5Sj
7DAXje+7Dw7+GvBvjv3ycRHyqdphG3W5xVl01kmS6fWGaa0Rjeyo9MfdCFyIqyHexKsNx03Te2Pk
Tze3EER9iQYZJ5hhdpkCauTzh54mpK1vyZMnCXBADOQVANvSvoz9kHADz15AEeDHwuPCcNhmtcQm
N2gvG9hd4Oswi3p6eMnV3PGSnIqPD0Ko2Y+FFGq8GplXbvtVRyQ1vaVB4QIyOKMdwRT9cpLomWov
FDTwHBL0+csJYIex2Gbp6MX3wHzx6E07PpMgyTNenDe+eKVLh5Eatc9OmigwK3EDvIuCI5bsvQ9E
BPi3uXCxJKVBWHYTsKJq3m0ZfrAdfOBakvuaYzfW163W6JvPiVfbvMmSAF3o1fPpLPl4PH1fTl+L
EM+w3wYcHSt5qXq/IWQ3aYM0m6bNI5d9goCd2hfrwXvMzbNxZG9RDGd7c7GLeJUJM9kgfaPErKkz
j/zx9HxdinizdsMrZomHSXtwdR44Gki4iKW9B075ooe+WoEkDaHzJb+yaX33S1lrTju+Cdd1EcYq
aatRSqu7t+rmoNylXdiRGNCIiiyoughG/vbwJW3Cx7bZrJLM3RyIP4d3NllR0cIFw5Qi/NnnnnUh
mRxRFf5MGuiOp/l3z1JVvYJIhvaaC8wMhThEZwFkSNNQRT7ijYi9RAk/fSRmYXcQ5W5JZbVbAWav
QuWcH0HlSBJUuiegZ5Vq0m+4AQGXAEGCEYGR0PtBa2SH5APq7Kdo+3gjnX+kOnm4TuU3kRn+Btti
g4beGA+LojQe3ZBOHf8kDP9vHHOFTegr8VOBLWJQqeuUnm4S6fq2IjDf7xX84RfsHmcvX1ItJLE5
r5fnY+6yhOQSUAiCiueMb5iooafLlN2YVPlXG5IZMKnUuimeo1+skPJ4V5W5bI2NcFQTofNLJpHa
xJvI4c4xZimh/sEV4/Gl7ZrR6dNPgw9qnfUFD00gkzbydvD1vujJ9dVrWTPK2okZLQiBSFZRFDXL
CdAKTURds1swl2LRf1BmPb+rzSPqGoUHctQu48nDfFrA9DS1QYqmzm7UJTRxRrztdFhjsanHpVsP
9eHxaC0nX9g4+RreodR2sBUetk0tJluji4zpr31V9AAtW+Sz029lmR3FGPrJNmLXhAK6jcZVIKli
OqEXZa8j7MT2po6RLDSjTCE8UzKueljCwHWnZLKYm5yvAaMH1WqNTr3J6kzbK+PSzSKvaZYbvpXK
S4slGw3Kkpd9wT+FsxOMME3WEy6gInmkgFDiz2i+voZOtY5yG6sQVD9F9PGlrNzJt6MC7OPs4H+W
JiM28GKa+85GIrno6TKjX5mAXCqEN6ITV5C6bZk95j7d5OhBgMfpguoZOMyXGipzjhcEPZo+KSrN
ZTZB2gU+MYX6/7SNxpNJ/I0lEyRI7laBc8cdMTB2kLASZvZ1mChe2W7lKJFp8TQWDlWydLB2TUJY
aEBy8gRKI8A52jf662oWVxdf+UadCN6g6/YsJLMdk/EBUB67OxbaQ7lN+h3Qxk9f9CeY4zO4AWr/
/+eFAS8lekY2oid5fFB8ZLEnED0KGPDbH+u0QexE2Q3tYDPy5EB8M14h+vJgXxB0SdkU2rAStFPr
gQp7y2u6XYpF7kCQ6FehbPkKPvPzZ0iRdqxLspNG1E3ANrw9NnoFQh8VOG+LryPJ/p3Vq87Rdkzz
9Vfa5W8hZ96wL9dLjoaoEgCkZsVkFzUaavs+UCDwzcRNCuvq4Wluiis2ymY80y8jLTlFSG6wakBW
oto19hcO7psFIZQA0xG5dsdFZBYuiGP+UCX9lO5vuVNcGIHGkG0kWovziUvmQcNl5K3L/fgwt7+2
TKqSfqDfKwM3NXqSXXyBfai/ilI6NgGFfR3HV2j4E8uzVvWBMUYRLayjfj33fx5eESrD/pCtPiLu
Y8lvJwHtmmI2EUft22zPmclObQxZKV5cb48lQRkOD6ZVmj4Jw8Q8q1OWXfwAbbDMMulbsZ/2iqV8
hc8uyO4wfIcTj56BJAkdNXbvNEGV6BRpbnPgKvopsS6lYgPdPnixveGg6vC4uWvRN00axshQkn6T
Amku/x8+ZZ0kl6ofkm82JlERZY/GiygmDW+szKTAu7KhsDWk8qjRMs/PMDRpEoCUBqqeLUiqSCKF
US3M4m0ZCLEmCcVu3ja3h5pP8eOz3ZRg4hocOxdtvwCgOf2EdJo+iyKXVSCjQ9KTz/DTuCGNmosO
fFq/8s8uboSnl+IVp2oH9dYrPHKDICtI50Us08i1YzOEZaM+Ms1M+w+w9zlbvDpPEUlfoskyX8oU
sMwAWt3Nn9kQcurtGmod3D0utph0yoptht0esIBzPV7liLRHclEawk1tX29aefZAs3sUxiqt0exL
qdYZsU05hAVeXtmfmcuImvTy7L1onjEsaCz2nq9iXLvLzcIEz+ao+AzbXiW3SNRa9QYcFskdlMpt
yImx3j8h1f60wbii8cjrR3sx2Jr9k5E8Qrbnq994bJhVMdVRVDOF2cAyflX2Cqem/6uReNzOD7xY
FSS2zzwtPmU+AZWx89jFsk6/XgDmCZxUC6y8AoUopYbW62j9uUpwcL1vn8ULENKoZf4IdzaFcfBP
VtpB7aN5t/xMCN2Qb1E9963BcHTFyrXYyxDh8jiy6Az0fnv8rPEf1eU8/EE1VzJbbQwkWg8Otqeg
AScxeNECgj/oJT1Sj+4ztP3uCJO+2SVSLV//OzxA/Wucu6l6djsN29U5FTbt0nmJvDy+ljm2mFYn
n8wv55Gk5+qzFSnFc1AVEfw/Mqw2rna1IG+T9KxPOMVZ0iuLtysFYnb3Z22GA6gbphqUocZy6mGS
dJu/XzRZW+qin4+Ph/wJvXAHDXKtLUhdyjUvepP5mFevP6Y2W2nNV1T8isHrDGucX0Zgyy/m4zNC
em12m2eS1LEeu3QISSXK24LF/tWgqZ87UwPzJrCfSQNeTqhpIcdHnOkGUYQj1ycHvKz07dbkLpv1
LJmtAjMOCHIu+xFrq1n0Fay1iFCUOwb7tht2bKAK1tkxtshFw60EjAD1igxK6zRDqGLCZkxqJD7X
uTb++/TY2qSY270ZbFSJT5MMWMAhmNUK7RrGn+xxbmNRyYCDQRMU4igwMN0E4J0HG53k40Dl7Aa9
iaAr8PvVYGB+wsNr1yJkX3N9Q47KptkVYaVrneAVUPd/fOMpEJ7jnJuJBMXENU8v7tC7P5d7/0HT
QMQTAE1nZOjA0urb1zZla+AufXvpmWaIRjYUhnR3cVy5DiAdNMtxJerhxcgIpAfndxl/5uMiLY5u
UQC8KbrHhXj1Dsv1xCkuC8Hyfw5GhgI23Jfdagf/i2jVrT8Q9d9i2QsQQmGz3u4mMEfV7xSAE6Em
923IJwflksdhZ5lCyIF/d0K7k85qKg4njJNmfR/kXLICOrsmPlqdKHtLsNSwMni/fbMwWh/UMvF8
LOg8XufB6qry+PiOuuO7PYe/yxnHNkiyORXkO+yxSkFbXtq1L+6zwy2YqG25TPWmnPQvclt2Chjl
+ISOoFMUoQRFprXMRJoywiSIhYANM8581TrnrZMKyLhKt4S4+jEzPJlsZibTX7yC9e6gwOVg8R/K
Y80YCT5VK0/VRE8ovxVc3qMEthbwdBYMxrVOGcDVuil+lI/5dnLWH1xY1VSaVxKFDntMScssn4xR
LqKFli8KK0excg/vOWoJ0zL7uKDV8FBEyv+HGwZAgvTRunXASi1J5VOhk1c5tMqcIDP+ESJGIbRE
F91bCBh3li2/Er5Y58cMDI6zJS/vD22/peyHPEy5p97ggaDXDS1o4A/0yuIfkrdVeuiXBjRKX6i+
zWLirMGKd6BRAo28MWJFkN6Pf7JjdBDJTo34qn3ZC6DuxS8jX+Qq8FL0gWJsRdnRP5i8LcMMbJbf
+HS1hB6z4aTJcjBnuEb84T6bWcgY63Pmvp0Gsk7xtoA1kd/JW/K0JtBKNrMEJ2crh5omc0CbHFz1
YC4Na0nbWZwqjs4J6LtBIJJSl9Taa/hglihm+p58fIi+ea+pAM0kqqHs/D8GRiy3fCdUXu6PEHZ9
MUgjUnvlaLsD+/yxeXe5VBAzJsCSGG0V6g4MLv8QjY4Aut3HO+hQdIvMCdgYxwXZou+TxVNdXC3Q
OKxZpa3lvK0n0VnsTHJfnigJQq2Dqr0AqELU/5vDdMShGhQvZ62JaOO5zQThAyUfU7XcYgDqCivA
FcxMUl5QydESEGxLG5VMofBig0qKvupTH61DBv6eh1fLpQ4ViIArNZcTKPc3Zf935J2GIbLNnEo2
mn8tnX3unucY5LoSj5vg0HaxZyUlLz4z4z+uv0tY8eSF9jkao4YCzK+gjHcHZixL5HFRyoXgGxPo
SjLlTf43+dW5UPJnV5H14pTTmBbWH0XtOojxk/BgJ+G6tgQngex309ZqmDfCZ/Ic533GwRbFJWpw
sAd9VpPJkjygaqyUnZ99WWCnXukK9eFRiEalnAmu1m1btrHuKNuXSEoj8fhQqKWZ9EXUV840J7aY
3eHLDuLajfMmA0BmcdBF9ZrFq/ELAP1EH06J9Up/cNfGIHQy/dQ3AjfVEjxaS/1xJXb+zUxeZuy1
LjEG1VIn4pPh3cac6SnlSoxwSUORl1Lr29r8G/IGRKWEyIuTBoFOk3yBjLTxZSpj/6BBkZAssnYk
E+fer/9uL+SImImCoymKTRdc1U8hhx5cvgZd1nQ9erMxpFK+9aTF5VuyzNrTIHDqgxgY+OjebB7g
ZTAG2R3aFu1baLk2cvoy3XGQOCKuofCa/nmTSDwm+5TiaeOLpNjn2Td02q4c8+hH2RHyiRe773r+
ElTwS3WLzUCG3+ro6CkzJ/0YiroM/WPjlYz4CZS1RMzC1XkNyNarkx/Aou1q5t1/zz1hWtmMeqrw
O4/g7tkRMwyCizD6QsdLTKluYRQwX9DJM8EI6XB3v6jRDWIGBO41nX/oWQCQSYTmvcUvx2xmyT8G
frv4igc5NW8dEQEzIZ7Im/RgnWQ0Fo82pmm2b3Pgo3XmKhbdjvYjAK8VelFvOIxixUVT6ISKWRGU
+JoLO0MSApXM1FAkBsZLkhmqoqUIcZkmbDw/JhPOdJkWKDUnaLMQ3IvCIdPRJtZLPzwBJEDPjh4t
XvjXk/VGmaHEOH7U5GCk3f2MNPRCpCt5BvCIK4ASAa7niMmYjowLHF0MzeIrvePrun0QCub2nO4r
HUA8rI50LyPbD1bZN2sNbtENiixRC2OSWDvMN2baE6pZJujCOspSc2tewhUas5tyG967Y5KYsEwR
LZhmKhUoywfNLAGwNmunySDKeEvnYdxcRpJ+wgdV+64JIV2fu2e0jHaljzTAqtYbJKq7+2m9w4pl
07Z/lha6MMtz7xj3ozZ3MFnEe+Sg4ZF8mrW5bwKU32TIlJ0VsRAxizAkZdEyuxHgYn6MEkPDqTAO
AHuxtJac5I74eMXP5N2OJCsDRf44xck6N4ws3ZOXvFy1cb3zgOkTPUdIGlt1s2uyUgMUBMmGbE2V
uFMaTh9ae7zoJ0LmUFsZVLA/CxYNAjWzBHk7n3TriTTsv0P0Lf8G2SVlau3H+Cj8ioXak3cDLSeM
jxnooFvYbj0TNmzIoWMeF+x/2GBsPQHuZccwuJx+9/lVU3sNpD2IOxDyAeZQeCbXwW6PQ1KbdtVy
8wGufGQXUQ1nwcOhyR0YW+7P8KSJpe7+QHWFy6uCDwX6G/WEYMDWI5BINQ0regqjyd6eCcD1rjpR
JlvMDkqlYHNGgb1e2a90p21l92f0J+CC2O7YF2wXJbgoVSVvqPOfdJSPw3DddBAm4O2HtdT/W6i3
swDPMuDd++36z63IkHKT22WA/jXExbFA8fcb1yTmQHce5clLRp9yCU1/0xGM2WoqHEs9yFwQfQiw
mGzK5D2zMk/E6fzaJvSsk7pFFBVm8vH6ezGr+9QACChVGR8SukQKqtZRVmy6V9Mpl02L3ClOkYEE
bgfMxkbvNQ+OvIVQ+Wk2rA2MwnXni4PoPkNql8dWGRCo3eJkvomR2Rq18BgcwR74vfg+zC0SKAkI
n6xK504+m7wYX7LcbiQ93ByVfPARG4PosSum32484z3WjEirY6GNl5w7EjIB99ksgZperkbNNVmy
nns1kXsApEgLDAXYqe8oR87LH0eho7RQZ+RAX+TCMcovrvlAlxGjhTwsIwAW47aqg2F+HDy7sxAs
+TZSi+sfs6BZgwvXuCMZ+wzSN0UKmaiOimkV7y6MH5lRHaqoOPbEkGx5Be/UHsthDnkYY868/TdS
MNRHeaEXdvyWizVIeOfNVCI8X1c+RV9uUlcaY/6I6RwSPRveW5pBLyvA5OCoEcu9to9ZfGpUc54B
2LfJ/GMJpYdGLcJleduz6oLnyRzGY1TBoOVxgyFV5tJDg3/Y0f0RHcdEUwrLnNP2qwriOS8/us52
9mf6BQ1dUum8yMn0ku4s//cMuWzpJSt+4f7prTAdeJKgWn/W4OEYIIuV4Dm2xuAElfKMw3FvODvS
3Y7mqBLZb4eUsE9xp28Fr0mnQO076DUbN23JVn4d/huOAl8720ixCEp60+qDFUCdd6F4eAXC3mhE
IBgr3V83ST6CAQbH+PDsgxDmP/xbsr7yUI1O6XtbDbxRsYNJu7h32MpIurPZb8u+sTEZaq0J7KY+
+bNuHhU4mEwE1GtRtXimE8rp/r65BQPbG9Gxn+P0QKZycmiO7jX613QvhbmFE3aTw8gNFiTGTs3y
LO5n6Kc1sfynKcgT9dD8ly99nkC+AA4TlG4ggiSIb5D2u3D+qTKunkbsQYOwhFc11sTw+c3RQ0yJ
bdw3umLp41jLupOvxvU7blr1dRSutsWjwRsyOJ2X+YkgRgjQl06VCQobXfJWCNyIX675hLwi/iaP
EBj68mCjuO93d36jrfWw9KVKxOq/ihvv8rvBXLzJblekRr4wYCuJtlFjgFu5rHe6qarUAOmm4UgD
jEsFLuE7HAB+22XcYtGg94ecEPClv1M8DciLUTcD0zh7QSgKTDBABXhM6MjjnHtxly545BgBHke5
6Pxczs/ZdU5Vyy9XP8lPB9Thn9QxOFFEi9dU+r36t2rrXBLP3ATUz/2VxqaxpQy5QrmKYxVA+136
exPQbVw0ManM+S4ENbYkb+k7AKeInTAesMw5Ku0yzVq6oEcT6HffvpwQvftD4sYfcUa3EcUNpt0+
pGdFEkeLIHBhcB65c2Bnyb/d2j3xuEeod4DP8nl+ql8WLQPY8KWXZSoyiCSLICZulWahW4M+mtRx
Hui0A+kWe4eHve1cZbSu6BbsX7qmU1WxfX6GVQYizn/LGBbE4jSEEM8pT6bAsrMPhuF3fP1OomE2
IinmebFHt0dKGC5xU6mrKqjJJntp4QvT/0gIqX4Rs2juX9PVw/d3fezZq4VG1yXkSeOIooUzC60W
qMg8jUa6r+ASQ0KB44rSM3AkXc/0l45Z5AvZinQDJyDI1YPGLurdvuGU7Vm9xC/ZD9SY4MopUtr1
VsNI5HVXkdvMNi8+mbg76MjcBlxbfdFXvcXIAzz7/ayOo9P1T97wwhOMCAMECiiel+DOi1Ag2uNM
kPgfkt/cfX+rRob4EQViFnKpqQLZ0x/JLBeV1QNuM65kWKwKrtFRE/B3XRTjY4QD5epMd5ZeGtg9
r0GONXq2LaydRdFJaWEHQ4hNW46C+4Asifn3PED/dp76hictwgxKxKWIeQY7+51Eq9gfKb57SDAq
uqT1H3A9CTThG89aLGfiHeRZaboM6TyioH/i9nlEBr17FUyX9ys0FvvdZ580FK2s411zu7DyOGDS
UqcWXbCvW0/o7KjvdSeIjnYjjqoptBJRGTuBEBF7pm2UGkkbBwwLF+ygUpBgoejHYgr3bxKPjHgB
0oBDfsmGl2QoXc/vTtuFbuf6U2HbpfjOVXDiQcM4KrWTIFxbd8qyDgtZMB85KEReQZ3RMNWVC9wF
XtEQgH0fgXk0A1ts+I/cASASqHESo6TY5bNnGWCltid+wGumOeUcw3+AsH537KapucmJL/L2y9st
Y0OkYGnRZQFvtAEkVBcitJu/lyINDGmygre42EjbwgfZej68pQTcyDjijcUH2lSJY5/6afMLObY2
0tkOnISN6Ge4pKI3nwL6sOjmdMt6CBY98APSRB36qdG6vUCabSqVD57kxLk2drMCFF9Vu7vR2Onp
BLXg95XXmz0C0gl8RVpHUxZmrIO86WqJcsk+2qXweH1EYhc/qX8wphJExg4Yv31M1MscxLXvzmHG
kIHz1VbrbfK0sQNdOQ0umv6jASXwf5T/GQio7r0KFJrOXvYk0NWh07So400ZHQuxFyzfgSeDvo+e
jdaPPzZ68J2L6SQIQ2oiCk0eBm5aDuCtu5MkioG7lGZphTshGHpl/0onQUxNBzTrdROr103TyHYn
KSHlGRtFlUFSlCf8stNXS6YuAndowo5hYQuB4WmGvMWMU1CsPvdsVVK7xjSBCbETTUR50ETGaVPy
auXA7xp8s0N8f9HZT4t6wfjSo6JciE+vbtRzHHq8jUHckUQ3N+XaOiNfboA5RQ1GDMCQ6Ne2UDN3
QiBdE2OSjijgky8onzNXOQcQAhYenJr9uEfK/rSVjvlmJG1JPuuWrZegHDsN+JSEZC+iSzc4oXnD
b0IrhVxOe0H/960hbCpKTK7SmdX4UGyBhLXsAEFRWxTCj2fYePLja4UkevM0QE44E6EQo28wsZn4
gAi+G1/VHnRQhby3kwN76fsVcsqSsU/lI0HvDZLE2V0nNvaKG4JinV/MHnjR0yRsMJVheoVEXq86
pqMhNYxfnwNO05RyYKwCSUHCXVTi1jBk+fVGo7VxfJBYqgXrtI9JI9vMy6agwygkn+stTzpsBX4f
MpSSADE63h7xgQ20v2iasEQgIH58I+UnANvQ7B/45xa6wEcG+jk9w0ZAVVDwxD61kjzibVf/80GA
TTQYH2SYLBXaUp/89AFAieliCeiD3q2vpfj77ruolp2l2hiemrwxDbTlu3YSWXXNqFUCz8M203NO
5P4HYZppVBBM5/h0NEgXY9OuwLKHJBahAk2dKIOFcZxreNwN0CQNXv55oxFicucGIrGLpbgOX/Kn
YR8VRQ7Xl19TOVQNurdT/FXnKpYg+mmTPe99TyX4hJn+4DD7TbCmuJjSuGVFrp4n55S/0RGDke6M
uIbPTi/EChRKBEB5jI2X+M04AIpBLUARab9xYmdt6B6woYhuy6FB24E1MgH3Fk5UU/jcGhBVYJ0F
Se4w1mmsNFb7c3tGyRXBWz48B1EeaGcz7AP+92Gg/i0B7ZEYv7WGj2Fm7lACqlKFmHw8b0vevY03
OkVV9b4/d6QnBVgs8zO2CndbzQPGyNJugZn9ajAA6c/nu9koEtto+nelcrhNjMxILuqceHX8863z
N+TErGmUeeTEnxmkJD+VnODnc0nDJJTgcxoceTzkqeigZzkSK89iOVW//QWCi1gd6zyTpAsNRWTJ
ORVkUyGS/7zKS33ZHia8f+Efb9usLrqZzBepgCgGvT2O360XyMKlWFDqt0AKXOZTgEiBV4WEHnUq
shLtcrXDBbkX8tlJ2+d2nZtiVUCqmUtYkkKCblcpWk7xMPR10zOGfaSoDuy78u4/1aQexIuViDpL
lAvFjjYIsBwhgbxnHJM7nIAaO5kv6OKktuUtgZz/pv8p3lEfeljUYbrx2pi356LbZuusq5FHfcxR
lBVSNzzbCn0S9pyNMQzHJwr34a3H2BSZwgO/x1c6/pYFbsxNmlkF4z/MLGW4sGF2/rVIuqtjY+f0
Aet+K7KxqTL4jHis0qvDRuks2gjLYS6NLr+eB9Po6MsbnY9rSHkBZXxwAofQi/5sSYadm7bc61uH
kiDm/PmEAGGJUXkapZVHIe8sR0XgWzYjlJd0s9WSYxnqPX5SbCzvoB0zSto4mzRj/UWbRRMGdNnN
1eLvra1ZEadBgt4ykQ+V7YEgrcJ6rmXy92aGMXl6eiilYkbCCWdLsxK22JKRfRhvlnt5FklHUqhR
4xT394/ijLzDF4386iwD1rkbJsklsRbibuJoJpC7LJsiigfw8WWKf3CjZvUf1tV1BxmrDb+XjN5J
5GyJaDtboDOiWbkU4bde6uDSz9trbSj8KGtj0GWosXz40bsRGeknrUaTKdYF71bY4OJY7mb0GMKF
BPcR23kSnRO63HliUqF4iLpwRP/Dt3wG7OSaavx/bHvvCxpnPd89umfBO599DqKnNDx5VSarVo7J
0rfbGiCa4QUPd0peLjK35mZ5+DE3nt9bZOxm7ckvRBlmyt8Cw68+x/TyETFWWBFTNm3rUiAYe5Ko
TAEe+hQIcs807m1pvzYhVDpUsKZpCRTcI3Srnm1LZKwcItLO/pSYr8JeOlJfJ9IpPBXiYaaKaTXE
/s1GLTzlGQtmYF3YK8IyTyZGuOKcE1e/WY5jeMz6esv0/rpY/qZGcVVaa2eisJQgG+9Av2CDzevy
Cl4+hFYkm4ncf3X7lKOSWK1y1eGQSzrN/BF3+/5iNN2t9GMPkb1ma4TydQEHd62/Nuxi9aKQDw4x
soCjijuH+ZBT9V9xrQzT1Y9guY6HERSkzNOwxYWmvGNPd2Oe2WIWegZzYRaQxtLpDRDkdtZTXw10
NqgyArEgwOZ9zXWe4nt9kq7+sUxLPyFfAXo7fvALAj1JZUH5SBZQL7GEkx9hplWJUGNqeGAq9YAb
zuC6qYOcJMPyrp7nmeshp1uM8miOPUIn4LOTBY3emr5yZW2ZMdonO2abqYsfj4lZrF7pbyhgxW4c
ZEoKEL//VjDJbh1EomekEna+kyCKckKdUj13wE+oixfVin+0ZpnOBLaC5v11GDhM+VL8SH5tuu8C
zvZ3ZQtBJr7cliXZ0ZpWySjOqh0hyj+pHK1PwMTdk/1eY0Ndk7pA3L8avOJ6LoQ7t7Fc1kKwV6ul
/hOzT696hwpZZ3WPVKMiQG89ni4J+1xj/Jmv5yHedBdRDPe7fOjy+xFTYV96ckt3ZN5NL13HgbFC
XM9YFnTNhvWobqjgWPLXyyINyhbErg68Vce7yxOEHBkw1Tz7HXCwQ35F20/S2B4t6RWdXeJZfcCu
6NBy8OfD/fU1NX5uj2u1zzVXN/Lds7Mxy4Mx1+RgElxbP1E2RJtYpItYAivXk+MJqs1oW7rRFsZo
1qhOogqovZds+wCjmphUy2KNMhy5IgUbZv5/fOjmY7sT7rOnHkiMUPoUhCBs5cD7uzF2fSz2QPZz
0eTvY+LVYneQQFr2pGY2IwShKbxgRL22dVT9okNfoL6xulD65djKTVYyNP2MevNcVBbfog+hM0c7
Wy24uaf4mRo4+JG5Czn5vHttycCKztBu8Gw/PaWV3rd3+mdyD9jtHfFxqnK3KwuqujzYmLSycxXB
vSK+Xb5GM46PPjXZu3QWbXaraq+nNKPDXWHEF8qrLjhJOjO3uh0DSwj4NQScAQmglTF0ILTPuwCL
lqKf4MvKrjzjgTBkMrSIu0N/JDfIqfVJ6mXnE7SY37Q/X07Tjs7YR3CTlVQ09hakYQI/ZOanDzqQ
ajFUyblLdfe8auQFEGIvUW8BIGiWMWhY1EPFIUwzcPgXNZ8p24QjFQYpmeEQYR7deBLCdp/L+M+C
ceJ6EG31tg4ajoJp3kO8aoXyLYf0kHL+xTCvfzP6ZuTnPFOgC2EP6Zr1WNQXPqDovyY4+xcY+d5t
OiA2z43PEFLHRXtfXSUhzb7Wl18zQI51E3mqW32dFrwvg36SDAoK6LyqlAbHA/VZWY8/X7OovQ4j
WgkiXLvgnPtVtuDvaeesuNbLDy/4nM5SUscUzONal6c6RqwIjO9AZmBnjuc3bwRytEQ7bqckYxpd
EhNmd/cWZsQUgTLg9iCyxmUZ7VoSs/POhK5Wiu4CWfQ7ldvcjlOdrB5UlXQfYyrDLoGoP2xHKkcq
jC/lAjH1y7Ufn7M/PimD6KAAs/4pgP6fAspnhFYm1Wrp1wj6K1kQgDEM7fMxlbKGf9WJnn3AgnMT
+oK0g9DUnnxaHiQlHtaMpyPCYyrJl4at+fS8Cv7IKH0ajI7p0LEZ51u0gTkq7zhct2BPLamg47gW
ZRcutJ80PD4x1Kc7LC9ThBMqPWtk5FsZtr01WRnh/yhZ0qBkypZfYnle482WWkIX03t8qmjUctdW
81GHpp5jAlWfxVJu0v2iHMQPy4LRCzP4THdXHrUZA9qz3bZdpcTlCvxzqR9bTm5onXaEpFmEf5Ye
eTCJ7JuDsrA0XpamLY/am9ampfiUntd/jK/0NRf2dZZWVzKsyaSt/Ne6EXI+LDdDJ/YGJ9pXRfpm
UwTKctyi1fAsm4l/w+Po2/Lvwf8b0PxLfiyE3TTnvqrmPZClJ8R2dghpIAeZtk2SVM6BEdenHe4/
YqwWhr9x2k/ZiL61ysWiWGk9tnK1uEHtM9KM1WPG2g7SvhnM36giDPtQMp5PzTuz/41fAjRvhSt/
wwHE1W/ALRyu0LkxtmBqWAqoBZdw+AgzsvrOIfl06+N/MD9SlDXYXuB+/SRZktwswWKYBqcsZ13J
vnoLd85fbnUdGWVRYkXPWwkbd0RueXp8cjLDKep7JUoYQghTdO90zEGdwloA9YhDWVCvN0BCVHaC
nZiiQQUATNt42p9idh+KjVyIlL8FOdg3ox4h40RarJiDhKf0W4H0BJLJskr/+m5JLSSp4mYiDtfd
LhgejAyWKlHvma2y8+dASBg6i415JzGe53hNheH4nTReGZQllIDO8EWCT03LjmH6HqhY+K7Sy7b6
kiRYFXZaE/UEIb9ONA35JSD+0GNQFFpy+m8s4Gxmh1igxaMYuMC1tfIeFJbQOKlYkyQwkMNUIm3j
SvH5F5L+e6VSZV0FcVqZK/EXuw2iXoScCxA/FJn8UK8xKjiJmQPdr5lDzo9U7jw0LlJjpJdXbvpu
lu9VbMTaXPk/RZI7lYQproWKRsOkgUbUt0/iOuQV+blCjKRmSnX3yrO5cURAMMY10fNgqqefwuDg
vVBbMSR+n1+SnoJ1g7fLg7ER3Fm5J4DxK0tjIwYRGZlKn2piDfm/iBHyF7Czxb43iDIJnOy/xlrM
NBpLc7Wsi5azoqR0q1FExhTGkda3hjO6CDSHmS79mmwrsCZiHNp6dF8bquymMDLmly5BH5oYR9FX
towLT7hbFFIPvld3alaz2VkQgObqzx9PbY/7XG+zZXVyQaQvmW6+f46clnMq/2owepBTqxLlyLbN
ebzkae37tx9asX7XSnkzQXV33o23iQ+O/ihksd7Vn8Si7n8XVFrdjQFU+1vd+VgG+Wm86BtCt7Zg
kL65LwJzIYd6255t+zHWSLKk++HJGnNsA0xLN/sOpQOhvPzqVDobxJTXz4VCAQdjBVm0lq3v/lL/
25BrILWtUOOiQ4ULziqC067eVTu62ugDaznddiaj/WuNIN2bym1givA6mkGYP9FgBwG95M+wl2P3
iF/NKZ2QCVNxgftz5GyGeUZ+54Ck6ZLkH6M4BiEsuJzbPS16EivcS7gCZ68lDOObUj0x53ZVwPY6
iH/JHZpKsWPkieyrD+MqygjQH6aTUqtuOQ0RYvDXy8a4FUF7Ztysdhp4+pgxiNrNTRyVT6bEgWLi
j/Gez9MfQ9EWUbU/x+wWEdfwn0mPe5lNpMoXvmW8W2Hiiboujei4gaigtaZ8zlE8E3qg8U8wB4Xe
qzH3qvvj8uA9N3VbirsCCO3267JlGm4hLxWBvrJ6hHq8s6L53MMg5Zt4dmMPslOYYdLQoO53IRlO
jYKSiCKGtAR41D69DrINp32x8H+xtZzSaemscSrwGgF9LEkAiZPKtVedRHpgFylN23uRAKkdpr+G
b0wRy0QIhHS74jeLxmSuuiqGvrUxzckW5UJekUgtvlt06raCgONAcCU8aAV8bSCQwCKo5BowUHVu
bH26ALFPeS/FRgqVpQmfYczpDT90ALebqW3/1Td9uShjotPEBryP/5XHl1J+WouUFGBrg/kohdA/
6bvjnFld1IEgc6e4ovB+gOW9ekv3trnPvv9T9zqE8mvpA5eM2xB9YWASjsPum1tEFLgA5dDxQYH+
zF7JgU28AY+9ifEkOuNN07j6pKsHVbBeig3Huv7BcEB317Pq6ghRUdDGrD9BAI4svysbyub7LY7w
aXTLo5XSXLbHPztlM4kVcnVHk3rC/S7JYU1JKHxng5f9Z8moTdp4P5Ss9essVhzTnRUiF1OwZ2Z6
toE++VTFhJnHBlR5WCVYQTOkRcgekZ/zhOOqOUfmASRbW3Fbk2TMuOFrDMlNpUfvug3tNEIW02KZ
gsn2udA2XKD4yYWdlYueAodFmFj6pDtWxmpB8ThES0+ZZwaCEHle5FedXDOag9MFWp1Pr2XuULDr
kQuDUrgrGYEpz8UEiIdg7g1T7sSKfgRxKDMHQAq8vCG6uX2dxkwu1MwVKrJnRk3R9sdeuyjhyPs6
k18hfGTxotjg0xWXKhW+qTcE7wnX/fMWhY8FHITmky9Uq4BhY1hRbj0Yw3QxGTLpiY8ep5yvQZgH
Ox7BkCEg0CsjtIiggFL7AA8NDBjGtwzqcwPPf8BnHbrRY6iKBOajYWAQ+rkwaidmoGjydXYLfSzi
b9dHcK7j1xsvOrmuDlQJQqAQ67j/dSp6POj1WNGQ4lmgJYSS/6FPLrEgaoJ48GEkPK8T7gJLb0PW
KyWsCdADzYsdJuIggf4r7XXt2JJOHR7VFN7Jws+hvAl6584tUCojMQMvb1K0SnlTlJPVOU+GY5rx
GFOG2WjxzDrVBif1lmAipIEbef+Yx+1xbl0BsKklJNkICBIqJH7Ui0SQswqR57/DroDK/1kBP2En
UCzPpFzDp8Why4ick9d8KCNPT4HfxENSo18Sc97uhWrK2e9jYQkw0etNYFzp7240ekgf4eJObXy3
zuJitBn3BMw+Xc2a13mPhxYwaY00eWtC402tcRuRbHjH5D283EIlZ3pNapPNIN8gL4EoLUcyyNsg
Xhq33LgYCXEgAGDFk7WVH0GEM1pvRMxGlT2JYs+0UDZt8Dk2+w7LALjNv/um5puhKqKJ764zkt6k
kwbFVPnhM06PXwyMgpAPehAUY5T+78BZJiJ2ukCfvksaFGX/Vb/lYUrxev/xmQKZUmQnzxehowJ/
Jlh/qOYKJtnmAJ3pmSDdPAcKAr6CnUY/kYtVaY5BfQeC/HDUOJr3091eZCyiGHKuSL3X5Y+YmGgL
jc56BUhS63KIGGBrYbtZ+7ylpsLZsFhEgiC7oG2a3GCej5SWQN9YRIJq5RfFVyE/7hIsNyttDaAH
OlGSlc6YFIqV7I1o19XTGRRS9kh5UtEhiXC0PCt6IK6gxibCBeW66ZA0mf7r/9yX4UanJtnaqTY1
3hRUQY6A5hIGyZ4Yb8r+Tu7+3xljgdo4UxT183r8/y3YAF1gXZKZuaAmcyI7Emabi2s+FCmqGg2i
Xs+WumTjCZ+L6V/44ytwUu6IHnbImpMrwXW/hr9cZFF1XGC+XPb99+PuHhqxYxqlUu6Xn3DdVKk7
yD6cgHCgZootTyFtwvkMb9aCdesYPLkOnYW1hyWgaqIn7JsYbodSx4T+RYQQpbd02eQbNbhdREY0
HuhjIdNOQkNwfL1keDgEMxFkQCFeGtSwsAQOJFJwndkLNzUTwRNobthK879/c8o+5vXq9zk4/oW/
eZqrd4a1BK2AbWpXmf2ARGTKurNswH142ur8+qdNhHOf720e8jO581BkjZ3DEZ1d6VJ0Ge6SbuN7
6qNWwvopb+yfD56mnmim7P38vETM2/CuIJr+bGrWWsylYe3awkCupmMZgXDO4mtblGWPpXMx0l9j
Dwfrh0NcdSQV+4kh1Uji54qCEVnM0n040n3GF26yEBkfTvaSvrz69QjC/jKCpmRTQznZtdFi1QEQ
JOi3YgMVUKSgJiz6UmubJ5rn6lVu82x8R+gjbb+1d3a2A3bYTDktbRACddG/nRbgmVMDb9pNLLMy
wpOUT/kJjxAEC4yAPd8BcmpzGtfhywC6W2sBiOg3qdvDWzMG4QMOgzQM8RnZzcpKdeTXfirU//zw
G6XWj9SigPkHkUFEr8X8NFxvMeN7NiYW46Lc1rvkemaSNUfgjJ+Dp4Nc+LBk1j8rSCk9/jxvZbUz
9JcxTWRaqOksHDRfj+e2o2omEI1lpmrzjXTjZSMIZw4aMKH9FMbdHTb7xQaVW1MLMSRP6QsoFX/E
1IZ9ed8VDeVAct7fwi9FPhI2fYv3hwsKMAyKs7JZ5IV0PMHiVosCBI2Q/0sxDQG54JWLR/WhaWiH
OjSdLpkgFGMdompwFP6eYx58Ii9E+KIj/P1a9IP/gGyGVnH3YJitT/s+e9ROxIdTZRxXFHPUjZOd
HQiynl6qS0Z/R2rh+Uut2qSyWtWMJt0lrITxsNAaqDl9qQT0HPvGmHLOWBNBamVCq9FV7W7Wuc5t
gfqd8Zc7Q4vRkGCCiG9pP1Q1gd8nNa6ybnMXSJWhP85ILEtHuF8Smn4Izjxcu31iJWp+FZwVGgQK
4JN3Io3souU8n8szbQIOq4o3dfNipX8yS/oQSvdssA4MbSLLYzI+DcnXFsrolduNLXdQbqQpiqAS
nCvUQG4vwdJmjLULpTlbKxpU/cnB9LNh5im0iCzmxTYpUNRYflO1qCIetj6aBq7nzkv5otTDmxgj
+yqQ4ol9oA3glhbM15isGGvgZPuqpBAqmaoJ7Kvyi+ekNSN0oVGdMW7X6uA2dM4FQ8q/h3CKrXAQ
zY2HW8+Z7L6igHksRyHiG0z8Hu5hji+wJnYXuDJcwlc3p7dAAiVY0b4IKjHUtl5Eh0qz6MUg0y+u
L42IZI2VR6AU/u/QSUWTHbl09wDM5F+QBgQLKKzKmXMKI0hfkW3w/yWZDY+X8P0X+PAGtIQ+sIDh
/nrWXLUIkW6EYj2kJ1+a/IMAbg5GDzcPGTbOdwGIzwY/uMb1pI9YH4Q7odgGrlpfSeJnwxMpXLEI
qGtJ2ah7LnJ+NuqJ5OYn5KORKCCtGvAAy9zJJeCBNfwV42hRQKr9JSzYbxWgy+6ajUWJXFDtn95U
rLCQ4U5fJin1Wen32KaXzkZAZGSf6ENwX5t2AoblOcPFLckJGkuY9smmJK2T+s6okVhN3zdHcD5S
TFZgKyYhubl0l0mMIXZCqLxdcgJyX0WvQUrLRH8ndRBK8RkA4Z6fnpauedfJ6r/sSXW5sp67nShY
bQP3ogN0+k/ENeVq+rwSV7ncyLR0VA27v1zJVhkrK9sGilWv5M2iBlZWVoboOhXAEL99LV3Vm3S9
DjU/2zLA+hHqQ/ZxTeQTxfZIeeAiMDp5U4PC6x2f34QX5EUIF+6NUYcJk+Hm9ZTUfYOJg1Z6983j
5uF7+dBOIovgeFCzNTml97eb4msN6oGfgcNnQWyD3S+/UMzJp3ZnN/HBGENQ7U3fjZuw07NMo/ep
ZQhMRY93/YItvE/fn4LoyzRbW5BmFkzpYLKkKF9QA5ebhyOznGjj74zipFwzBwnRtzfA7+q2QsIa
FpZejrDb2ehJVNGY+9vlIh5QiDcYKDdyeWRnhLnGENvPlq4QFnNrmdhZIVil68T7Oi3CW+TMpw5+
6PeIwATlSjCQ7M49AM9D6HQPhRtr/Egsk2bPoLTI//BOWA8m6h0dwBemq8gdrRIH/phIF6SPEcwy
1IQcFlsyHFgEMNum4yRelqeD3lNAVXI46wsUmKlakhMn55Otm/RaiOe91fEawxuKkYpai+tXMM7j
1AmUMlF7MNHcUjrKRCJT0z0MyFrQVOyY/pF7Tr0WD7OrNf60/m1AO7cNUJZTkBH4/b2kfapiMx/P
FK386wicPpAwG4lAqcxMwQBu4lJslLfkvTtpUbvaRXtRro4n/2LRb5JvmlrpXZm7pjL8KuZ12dqm
IZKVqEDSAhcV6MjFpX63++kEm/7cVApIr5pLV1O1AZtrCDRBmdY+13hNtSWED+1fE7f0czP9T5kG
3GrqmyNkXmHuUrOKOuVHsHs1R2dZaoWPn0G6aIXtmnQsZMOry8JaFNV4+Oj94yRW1/nu5a4AjPpW
Li9eqiPJ+fyhh4ly+uxO9nQJk4qGxoAJtAf/jAcOYXnzBsB+NPLZsUgmoOJ+fBNMWz6ZPp2+f0r3
HFVIdXpdFbgy3QqGsc320YOuT7DyQLZHnnF91bGXwvyRmxNvVT/VrWxeUGDKik6ZxlPXl3/ei6Nn
g7ym1o8bcgO0sZuSwsRzUImMgcycX3cDdDr6ZXaY/HbygbCLyDaZUIceJ1f+grJ44NULPYfwhq1c
oWCfjBk+i+pYI1NatnVIYJ+OZvgRhb0HAsjxoKqfMa0I+mXns5rIZz4SmXPkTW5Jm/B5R2RcCkRt
9u5HQP/EARHYcEGT76PGozp3gm4HcThWMCsLedKfzhcDFfmBk2QVEQ+B7u4Jp6Q15pod9xbH4/wB
JF0ltsEoZUG6ngsNJgwZ1TolaI8YGtfA1vhntm6onaBZkAr59xH4v1ptfa0MuDtif5by56abyTF9
us1JoV6qB01tpnbKuAh2CKnVKo4v7nK7quOnCVSx9qYhlzHBMPiu+E/lxyzYoylYqfdK9sQ+ZU94
EskTfXOEyALyqJyEI8sI2ztJCa3LGgVKRb+4KJ167+0eB/j4xlvi4vQLwerTHE7kJ6o1GC5q+QdW
5DISZFWzFsG8+YBIOFMCYlDFZ9FxZA/YfbDjSR3zp5+OapaqLcpXL7MGRqQ0LCRmFFf0yjdOMvKO
uxWRuTddeIBmPoSydCHbtqzKZjFSlH3gYdXMgCM/aROxa+PKkLtegaLNvLvmGGZBsvhqJR9DaGs8
N5hVkc6RpSTaieyeokpBeRq5fO80EeXLzylyfXPIkq2RpO/4kblDoUicgaV4eR07giRpZv2BZZIE
EQQ4gB1kpDLISYgDFq3umO8G7ElJRVqjENP0TZAy6QOS1FTGwzc6F/W0bhglQFIJVheHycPUR7+Y
HDpjciWZI8mA6g3o45uS+CFs4PoQhGK6jfjfNMi//gJE1U8vCOeGjhJYdfQvT32TcnjJBLt0KdNm
eXZv+NQO0jRvCWCDQIzL9810UNKAv1e9iA+baD3VFnFb0PKToyZKcL+7dUdatsvyuhmNmWtU+M/K
3n8vtE3xVOm9MLvKHRj086dHMxXEWNCANQfgPcaa+OK0dE9ZwSbQwKdLTnOSjp8UKRO2EsBgfrW5
WXSSkZnFYbjKgfjq2XiJcicm5BmAZwDlLu2BvGdAzRPWE4tSkqPjE2845KFue66kOuY1MhiMu6rP
HpsuFmaP5kC3NN0YiqjjoLEnwoWrqUpTpCF1mYeylSftbIqvZYKZAzbGndGx7xvVWlxyZfC2gOiE
G9rQEpT9wbknjmAwQXraIkKZH66NUClgPgQEgfh3gO5IWJ8d8HjsrkR2oX2teWMAbJWrzKOu3TX2
6FAoLIzm+f6r2q+um4Nxjdq3kBsgQlf18MQKHd5X6uZQvDfnlkSiN8tA29sqlitsvbc7QH6xUGDP
g4MYKSXgqUkNYmWxiJl5V0mX4cLaJ/mMmskrWmKA9rjdXDupUoiTd7LV0v6h2L54j32GelI3dRMC
5Kp0ux4XC0ZeZUZUgS2XEV0TH6wG7n9a+39RlJRXixuRjOkMj4VbOjZxEm6qw21lvP+ZoZik9xus
oHz/J+el/gugWoTFgVv9WJox/h6j8VAiM/oitKqEsYBqMZupKQT1mbm2f3RUF5l4nL6L6A7iune1
qSRHc1uB1jKEhuyJact8l33cIXR6lUeTimfbKIRkVoFsVXhOOBowKBKkYI9JbFaWKn5aaRfoy0WJ
0GkUcE+tKPz7lzXLKAvNsXE87YPVIAoacyeJkm7BsJNXDVrZc7JOxlDFJCOu+mpJIRVd3soDltoj
vDqA91B1vx62YUUh0OpP+kmHe4mf0+NICkkeQzz88x+hOp4q0AUaybf5nzx+hPU0+1i+bb2xwpYL
/5TeQ1ZDP2m5qJ+SbnVOTPzKDo3x4q4FzTYLpwHEehyYthT1EHm7VftXPAtPKT8AbvrJ1BO1Y8RX
EoHYtRkei14OWkMbuCNHN567DMG+x7j1YTHMpNdTfYiZeA0XCOVCg/YT/8vlkcuHMMzkKjYppP60
+GU48pWviu5+wV+WQP9o/wFhMRG1+YcVi5xcBQt+JEb1HJbUwNhTVZCSO2p7tFHPf+1AmxCAlWvA
0YyyPHHz4iO4tnrTgK/f2rDfDAb7Hd8Qh7ItxSfTv/NeyaWNS3mheL8Y5qOztyOcgdsLYyKT+1R8
f+veCP/OhjImqD26FcqcZUb31ZAMP+4+BECoLBuGZQmyhvGYflD/CTi7yTwNSlYLwKgUI73wEsSn
Lz0++2vpyBb/Do7tKCE3u8thEWIqXh42+ufZqmSJBfcHFFu7slZoYUoqrvXyS12/Hk+I/YFIc1aM
bF2VDJFpgxDe6+dsx0HNvMzBs5BPhDOSXnXRn26NMQRHF6Xo0sPd7BKAU5b7wSiXV44zX1SOLVjH
fN5Hk9HV7psGsLdqV18/V58KXd4wbn7ers+CIbaF1LyZMdt0D9gSX354gjVOJLRrQygTsYcj+Gsx
IFG5mrYxtWKWFhCXHmxOWkLx0vCvZnU8QaXZ5MD+A00MX4pR7I7bIIBRK97qHQuSCTStFHyCXEV4
w6jbTLOCNbLb6UAzco1YGFadyToPZKYBwq7YkmFq1mvgBieN1TNj0szW8cxKYBopRfkoSLHnqrA3
d0wtAseZj77KkRjHIjPRlkfH/qbV+8pZ3OR/dZUBCZPCKgjhW53SFj9dTBGVOspFCXhWi5CxXHEH
/HE2Ew38r3/Fh+APTeTKWONESVg7Bl19Aza0mQxfRHx1BlNqN38WXbhtrnPZP26w8lPQDP1cU70I
KDpQVwCJVw/r2NbrDPn1sT1k78uASPXjlDzHtOFQvHapmJw8utcmvS8TJsADmZev/H7G8v57RVe5
kAgztVhNqUzRH0JxRH1Al6O26bzwVX3+1qtyXHNZy3NGtuI2VINSk4L/w85b6/3jd5/6zgFUHTof
GggxRqfMPL5W7rW4vh+qxaSF3H6NySod4WAIK+yY6L8yFmS7zY3MFrNe12pZHA5lV6i/3VtUSr/Y
/42odin63kHwBssC9PEt8RjkuHJrumkf6e1pf+5SkeShgy35D+MdQZ9SYm+rRMX6K3uqQRjx+Vcd
LTrulm3TWuAK9njL6JvhUjTZgy90XgNWY6/l14x7H47b/axCJV69/uimnK1R3qsDF58j+rxE+mqf
G0Jmst+h7UiS3ZkRTwuMrL6Zdaw5/2ffvDdMtLiJUCOWEL7TYUhOirQVdI0lCSjFoCf5moBvwRjS
KGUjYd8pI7llAu1kNFbSrr1Lven0eGtKXyMPxuoYoBNx5bn5DbbCAONKdRp5sqzUXIFfB5OfxJjO
CN44gA1pX0VuGbXaOnyyUMEfKnHYDrmT1CjVGceyKFtdL55W7SmdtcxihAnyHjCYATxFQwKpBSRE
SjFhl27hZ29RBPooYl8nZvqyWxHmMvIz7F0oLobx8L7YHonW3n0soiCN2B4DcIrYL46H3ZTsJ+Bx
xRn5XuVQc+ltdtkhWWqvWADKW6mp59dDTqzcOBg1R/r7jE5PFHM7kJiid0VENbXWsnx+cKPQVSGx
64a6DTbcg9GKsFp25UGbSPXJV0w33XLN6BmqQAEBStyhqFP/hE5smnpkgf+VnE+4JJ0GBGh/Dapr
adQtaCULv+DWmZzlGm9y9Eih4PNqSEiI0aiAogrr0Ks6iGGbPJUYoBCg9bscS9fh4G4v+j4FipvG
EcOsXfouSwim0Xa3Wi70UQo8tI5bxL0aWhMRCM8W879vWvOLCfC1q0oM8yDAU6t0wU9ghmMpDvXx
U8qKI/QecTQKUdLSJx1er6OEqdjW29C8NmKn9ZcBFTJZIwItgXLcf/cc+TIPyGlWzfPXBMrT0IWA
6znMTAFMnUb1juzBtFRKSwG5qaqv2nU4cqOnYd9/yKqqYEeLhCkv8I6OgDiRDVOn4wswITt2aNK6
JObD0pe0pPwD/pK5KjRmBIY3ptVTmCFnEhfMiY0AsiXWNZtlty+DA4cCXfCUYBzzeyR1cC2BLS4h
/rRVP6y1YwYb0Oj0EV0RHCda3UABFNqLX0I7ygWdT1e4LW/Hn//+ueYQkL0vYb7xHsH3iF5EkwmW
U0EUvUjqqJWBQLik/JPPJk0AOKTAwRh69Bz+NM7Y6iPqRV7B58NuDrzMiTf0DqDMWxP6CXUvJCuN
nJP4VjLADWiTcs3R6WClWeU2mS1Ll06//40jjg16ZCM5qCtj6XIFORBKCp4OWZJsyc/LE6weQhWA
G9uoUO4r/CqM4MKoy/974CQVa5G+nMvhLAabeoZQ2e3BGs/ukT8Z+V0Vcrqc3cBUWOeAITFy/t8o
WD5YQnQrEs1kdzf0YmlxjXLRG385pJQO8VUrEspGPObfAAB8lJ3oWUhUszNOwuDLLpbxlEy7iFDi
4FaYh5mW5+cktrkhOUgPrnT3uua0GsukDPggWmxuaNigVLClgQWuhXRD2xllrAGP1D8Pfd/luypD
EI2OooSEgGLJaSftRmBPGq1mgAOx5xF6psVkoA3QLJwBwbQ/vNo/9AP2aN2xM6Cev+vpHGhsNsQ3
9Gk+zwPxVzqzd43GxFKmofmm2j3UVzDjtqGuU2sXA5Wl/M8zH/4w03PRhDCKf2v9kNHCUvqGksnT
/y2+wb6XtJy5F+p3DpaT6AGz97d9qBhkItjaTYm5eeXbR9kqs9mAiIgw6Z7jbCHtrNoKG0Dr1oeS
XSX8UYDE5pt0rm9Qs/x4XevmssEeOZ8So+ntEUa7kaJU7LGVYxuUs7CWN6hKBdvA0+vmMqMttJWe
IwwDKwPh7vpURJ9yeXeuzf0XsB1eZ6SLbPGsLS1Vsqbb5SHnGSKLdOdR1igYmg2CtH1tRseLygns
Q462Ob387JecrOxkfhJexJq732EwyvU22XCkG9b+DvQRHeSvD7jgRh29jTuC4q6knbOSD5Ow3GgC
R1jivgOmkEQDqiRlXJBLMOaEMasCiJpf4Nmt/c4fPq/hhMG+vAhN6Bd1GCscgCQ1MGd3EV4LQOcK
25LNYHxCJhwF35BzCDmi3fufIKkAwH1g9Rt7KJtVE4p+oiCb/1SgiYj8XHzO7POEuub9kMD0wudw
fHNPCEVx1M5TA9HWfqN4dfZmPrDYi5aO7H0V87216MBjtURDJCGCeh9IqR7dtGKwx7sewonMg/IY
B7waCNFPuL+5uOC5s6TMp122ugjOi9yTsREJsgnS2OtJtjLN4poAmNIGIKeuIGYF6P8RV9xiRjVD
uasohnPOWM7+RcgKe685goY7Ksg3ASkYKUuQ3A2wb+RNnMM8B5cH7I45l4M8kN8YuWeWDaAcA8WL
yIz6WEUGTfObvj9uqWMMzaYyaFrN4fNpEkAVQlZPceay8wxas/l4KGCJU+/E6WjWm/kNWhgxKkW0
+BnkCmvNc8pG9/vf5aL+K3h0BccMzWhGTmKfbn3erpkkYSiBgJiEv02Q+F+GzIb9Z38mli59mn2A
AvxIgAOzMJ5YsDGTeA6T88733f4/8w3Uh4/ufNHmEwjd0T3ngYuO0XK9Ik9DekguSaYbvbWp4Omu
LQzWjAdha8c3OJGWvB89M24Oini7R/L5E8d5AKBUbznf3b9nNjl0av9gE2bXVq1eYBo49hmS/QvN
3K+iSyzZZ4T8SlHoDhmvGeqDzuhag0ZrheaarfP+uNiCbhtRrx6WEkDkTZF6w1TjBuKKJxLrVmqL
qzFrwv4USXDtj4Th8rOiq33gYnLqH+gaMq6nxpPCuOLLpV1vp2WnvZJmO1L9Dp/LBmUcuxD+ivnx
b4mMQ5j+Gais7xDqwGURE57H7/YmZBOvQdab6JwvnUftN3yis+uc6eltVYktAa6rsn4NCUqXPfak
3NSzIQ2obZVxjXVsdIEE2o1WT50LuEoOZW+gSMA40LEZUMfjk5zGXXOBbXlc0sqdUlUT+tBM8Nzw
SoL6Jm0VkSgLV4o4MNszQea5xMP4YwX24GKE/jXFDQAxaTGv3ovor3OsHE/K178rR4dUva2jMKqm
9bakCItGlKlF0IHyK6cgKUumKvbUlFqiZKGIpBFrhN/0TmnqhYdO/EzhRJw4CZdz+8/7ZVP5g2JO
5IFyLAywoNmaoAyFw/N8LKL0jqBKSWmL1EswwNlTEvqFBFNzBffuvDszVQvvMpFI8KWvIdAvFVov
QCGCZ/XO39b3iBJbb6exMJAIvaYJHyTxSxF8R1Wtpfmafjk5p4bh/WY3xaXdckwsx6bxkI0ZkoD7
rYNs/ndv1zlKSZNBWHcoFzUtpJ6mXqdewb6XSTkoKMhFiAwv+f0xiUvg7Npl1Wa8soMdXfclvE1j
xb5Tx1xy/6Fnu1Ak3U+I9L4JsUlUkHsrqZ3Th0IPHmbgCs7kasA/iv+dUwPBaV+8pStKjQeVLVMn
M7g8bu++4ovMKb/a5dcCjZlVdJRCFu6zwGRZz6zYiPVYPfCqilkFnb/2z/Z7VQGIX2BdfdyACSzu
BjNvZfZCRY0o9XCYPKPHb8T8WDbYy3w+HK/0zDynaytoZnIVjrMwWBK63WicbX07XpBDATieFhHy
Ankk4Dk6gU+dX09ulCG8nlmzVMhKQOo1NMY6uUiVr5iF4o8tKkEcPZ1U4QFhuHVlyv/E91Lzyj4X
ZiuCSskGltwQ8MHWM6SjrL1oDBN4z7fkODecKYXU9pPlR4x5J4DTPI//DAoJUlEshswSzETHAO/M
EeddCtB3PtEH0yGCSd2EI9nU7EE1QfZ/bnjnk6bldzcV5bCBAx1yZK7/Xvgz2dSmmrpgIaCINWqz
qeMzmvLO9U8QSdZ0RmzkQShZXu78E+f41nyHlwQktCxWzDR4RtIhtgT3GSXxPp0UGAVRuqF6L8fw
5JqKUapU38vNclurT8bfvs/MYYEyF2kvWKyBtBr9hpXx6dXbm7oYWLpV2mhwEwP8CS0AT7eECCfC
OOMk+clVYupSpKBJHzW+dcwX3awC8OMwQqT7X2g7Z3Z4f6AN2G2XP9DmepyMq5ZFPaZDVuw/G98w
jKU5IliZO0c01HkqcAQSd9EBjbrtT9OYdnK3t6i2PH+CJ5UoHmSpP+lQVGgdz9W3pr9hPQmPTn5F
fmSARYlJwYs8sZR3etbJXSS8FMlblRgGF0zXpZOKU8FlTN9jAT2Aa5h6CJIvNJvtZuuJ8U4TzUnK
NyOveEpLI8yNkDE2aOqTYbAmMY10BaHrK1PP/vKeC+94PvrNE6BulJfG41Lv/2FCrJggTihRQHy5
hwEkYJvaZJlkFxGb223ervMkYGa2d5ElGnohLXSSBsOwmyopZgD3+7aiibqGCRksojbf6YI9sBW1
Y2IYOZMzVp9pS23VcLrQ+DPse91Fgy2ma0a+R8DbPJZ4vTrlr5OWTPVezuj/jjKBfg6lrjJSywFM
L0ol9+FDxP1sMrNpGKCyE/oVyGMRCGk76hIbtKVic81R7f2oeoiROP9REt3RDlPSQ/82jOc8Zvq1
hzRwyKHh6S+91l9piKiq1bKvTFfcPZ8JAJBfcg+g5xeLIg7ZpSqXJ2J1kemZlGI+r2MQUr0jz2fi
bqxcQHCfk47WBtVxlcSKskc68d74RSvaAWoe633NzF62DAQzrVWVydRT8HjQWhzR7Ar3BEXGB4ZQ
F9P/iZg2TnM9698faPbrrVAST+Lxf9aklCDd9WWHhEyQyI/Jjda41k3TcJ4y6pFX9hnRwUa8O+dU
lGcwaDYhWaor79hUcH4eZrclJhxvvxfnnrd3xfhOZZApHTsQ+KawrFNeNXX5Nl2OpLd9VNgFOZ05
ZpiLNSbM5D7dDkeDLFALFBE9NjEKg6FboH0oWpHTj0gsfgBCrQ0YAbqTtPmTFemB8RMGFBCBk10s
YtRWizD0vnkq/j7/RSJSr0qCZVwJnbj+XDiff/S3Sia77KZ3K62t3rrcgXexTYZB7lwoZ2lDkgRW
qyu+pXt/kS84MoRd32w4AMvmXESZJsSMuCUO2pW6rDzYRh9jwOCFrE2QZ8SH50RqbmlD+QfOvAbf
WizwPUBY+FTFiH6yQzxqubb9UZ9ccJ2+1hLP9YzGf0RaXO2Rb8yi4JK3iRu9ZB/H5N4yS5QGUXHD
1nDZnlyJNT1Lq3USVPeBH1QSUfh1F4zkSsb0Pc2ult9zX5MmLY5k7hzQoThAdiBLbwj197+OC04B
aG6ps/rHQ4u+rJp6ih/3pG8NNcNdQGwCuj3OJn9oVWU8cUzzj3zambo04CSJfDy/H0HvhtwX7r+O
i+HAbiJurpGrvp96LwdsxrL29kZ7tgaTJ3mWlq7XqKWWpdRGbaT096qYWHc560lGpTSlMI7QtxMa
MpkoczN5+NgKCzWI7Y3vEZbQgTetmnh3IDqsqPSVARotetR3sYMr+p1jITgNVAq2F1i0l3pDDRHM
CGk95S3TA+cgQylWjFRBSnprFPiS58ER8ijzB2Uc0ApNgJyIbhPxC4Znqn3ANEFaI0hqY0ZssKzZ
3a5FNpOaO/WYP38BmUtenbb4ttl+v1C042m7d2a90ze815sjFPMP/qEO9/Lm9ujbi592gtLmLFLU
U9eSBE2AO4DUDaAgTObMEj3VS/tZ9CbDMCcH2xZj/Zio4C/mtx9q8AVfga92jwjxoK+o9uvA9QIS
sY7MlW+bDWEcQMgGo+sqqClimywhcGqBecUl2gn55p5m0hPxLjpWfu5YoX4++u+xrHM+OrsjOByy
0bZkpLguRn0rJv1plcQ6uucUBAuAdKn8vUD8NJ5WXepq+aJRgR4hKIYJbhdkI7t8it5HZwd4DOFh
pIpvntdkcFz+/hTikJd7n62PaEfQ41yJqlioe+FMRVSWtP4eo8OLEcgENL9+hfkRlgCW/Y2rwFwR
pivka9aDGqW16zChFHpvJVEqCOK7Z7YdWlWW9fHffYi+BBfxTXVwQB1cLvCmT6bMfx7rjka+CnTS
CLnrXNi83yuzI5ifDET9CTWIDAEjjnwB8DyLkK2zjkWI2Du8bXniZEeRb4tSQKMA5AKLQyFA9Dwe
LpqMmjYQQRJSnk0Q4juEMsxMjUgPdUSrDigT33PXrEA2tNyz1jqp3QPNqy8BSGyMjAzRmV7jfZjt
/nDkVYzPeUv2FjSneGU68jREEQaXX/giyeT7NgROWYda0MgYPPFXVfT58CxHAf1v1+iR+/+Z0MUx
br52vd0F0LpY28urK0LwWD7B8WAhoogtbmVbq7qpT2HrFt4q/Wp8+6jOT6yJB/39HbFSi2AQgXBe
tmORLu/VV7a1g+VPjk+sd00J9UxXTeYwbzXwbUndp+hPct3qnqChp3BIep5tWUzeReLQ6YWMDTqm
64EXZ/twzEoL8wjIu0PHB2y4YjYKLx/PcgWuFOd8m5chblteVjRzbUolmvRnCzP59hOu579uUlOs
/CTk5Yr2Bao1/NtahU6baskSGTi+zqrRzCEJgQM2NW7LOnB38dQPqXfx6GjPt/zFAGRSTvvpRARg
IcQU5KeL0ZTxJC0fZrvBJE6QyVKhX5NFm6mwiJ/lP20OwibOzeBKMgNAS4u/VsDlN3LU7+V/goqd
9FeW5YVs22+G3PxPFh9MhyQF1dCX7Q1I813DNmAYWh9TdYT88OEOlfbirwQzcN4x3x2fjOq+bjwd
aoYjQ4rnAIsl38qMT+4zCcOT0n7sZMW2dIVa60VbWULN6tgpZZ755RSxznuUwN4P3exuFNU0noaH
cWfi+vXD5o+Wm1VCWlbC5UQ35YdygHZPKbPQ4LOJ0XMphS2eAksnkwDPHmmQ57GOo7YW+prgsEAQ
NpSRzGFZDO7yoj+pEHdNcaULTzCi3zxuuYEpOqMN8QIy11NqPMxEPYhRJQX0ezwSnTRSk0fWk/i5
6dmpVCgvd3DSCxt5LPcHSKi5GxhqI6f1xveZBtVQVrNtsH7V6tEMG3+RD4zMGvtzEWKBFsMvPbAN
SxWuEPQKukanwIWmcnjWUGzpRSB892sW2JAD/7P8m3TH3cbxKn8LuiNpveI9aCIEV9v5ZjkpG3eK
HMYRbMK7SnMIdWKWJm3Mhd/Ww939tjYdWYtqb5C8kDPgizk89+zxIUDmY5HO9X6gdtPZq9b3QqS1
iPbRO0lkyg+q1V2+vp0LsakbY20xzZDleX++ZB//FIMDx/s+i0ejnUAw2bE/0NlxSAFxd2lAIzBJ
gQCr/Hiikgg6P6KaL0OpCRlRGXlXC6C/eSulhFZ/Rt2r1kUVDiYr6y/7cXQAGDhjAcRhDUyzx6pP
8e/8re9fCmo+xw4c4oJx3JwMiDIVQG3xnG1R2AfbnI0BkLtd3Mf2rt+ZFdsZRmfJnaF72XlNrcmW
X8lzNJ4g6CgVK88TI1QoMEF3Yujg9PGoWOCuNixa2T/C6B8DSNj4j+nIKnKFfQArGzeq46RtSoAt
0TGd+8wWAFnGoF1+rD14pbVGyWbcK4ZAlsOMw6PX+9c0DoFt4rDTit6/RVaxlXc7r8OewqzS+vlU
L20uDK5b7ifXWrIpIe2dra9VR5jSYWdyV6nWIDqYH17ZsLoWKKSy147Q2sZ7uaNo9X4gv+f8iY0Y
5exqQw23tBnc1sEuTW0NxjQ2wG8hEX/fBWXoMG5prPL6XSQ/+fuiH4Hkv16lYQG/Y3xTDKzThlHX
X5LCFCl7ibgygWvNw/jtVvfmLAjQces0b8o0/XUsKkIiVkJlq3wJLJSAtf/9E1IZA4IHHsMIyJH/
seD4Y4mvcvvMt8P2Rab/Pl/HeH3/06MUEdtHmef1mWB3xANerlo6FLowvFfHiFRekkYiN8F8/SB9
mCnc/vVBohmtH2PfyCwlQ4m0j9YXkagDWzCtT1gCmBGDo0zBLudWjU9C7hr1ZytMErAszxAoivaZ
QefJea5QdbZel3i+u80k13vGboUnJJo5QUT9B74hIy4C1KmT3Ygr448bRwk7poGwinOl0Yd+oT+E
/gOk7YdoUoHNZCognInxl61aKIRynu+9uaqNEQhdRNSp8sRN/Acr2PnThFVz14Qfk/M3VtI+Y4eo
kqvfZdrMCnZnaiPHukYu4guFXlKLhJwZbXmW8T/KAY5HfT7l1mwpQ2jPJnSOyvMGfCwBEuDvtPSZ
9PTVip8QZJcXFbyRffvfbzIBfzblFmxmvocOGu2Zt41SiIi/qUpj4RFO9z5KXH4XWaW6uH7O9LZn
QtJwKQtrSAQ2+cO32Q+fRXpYZLGq0IYe4X89V2lIilmLGT0cYEf2KsL0r5zinb0kwxpJ0dHws2nr
XRsv0psN8Ttdk4J4AS8LjDhTB/1XJ+wm4aad7VtHDpPoEqj3OlCkcuK1ex40u3J4gbEUAZOb3C9u
NfjDO/8hfoBypwYcl7OfEVQO4lZlKLNBdEkur6LrNhVxXmxDgFsdCceamcZ7Xbc9jPxNQufbmduV
otJ05k9o9oZoV7PUMaz5SN6N9VffQ9eqiOOzFwNx7RczYnvZ8DuazztD0wd3VEAOlakKQVvozy5e
QDvIC7eeteLbkm+Zjyv/VzZUV2LPliUic2Uo1Rp+3W33AuiKhNwWdMHgq0PpZskz/KxaMHK0ikB/
EIhwc+5DvdT1ZtXvakYStjZbDxggZk1v2Zbj96/lZAG9QBgh2GDN/CV/eRWTdpjUm1i8NUVQLeEv
Za2yH0ZwR2FFZMorSKRTILxgSKiz/kwdDZKsM8MDqmUX5sgOrrzM+JTClwgttltxRFiI57VeAL0j
CoX8TuOR1d+Yk8jnSwMKc2gE4YEZ4PVh+nLQAXOXuYsu2+sBE4i6EJVV8eYFT0OowvsZdYhbdety
aL7GR75SWw9j9YcOOY2FJtK69OyLKveEsCJkSLZwfkTjCojFFNyug54LeU3fh3628+k4nwgafco5
rmo+N1C/5m6ImIGwLcwODS0jLNDBFH/+6KRMi6Xgm2P5YhWXyIV947wk8E0IwsF09pmJXEIzYE6r
mRNW0v90pKVdSMg4lXkc1FY0xtF5QrfXiMAG/8QEjqrL4OPoOHzSM+S1hc8bZUg0Ntkll9JjgBEi
hDttVSV067fuKjcdvVWQhcezPGkMRueukDrMhQPS+Hkfp0WiS7d4b+h5Ll0a8AC+m47ArnMXAvHB
HIZzp/L/OwEn+7kl10WUSKOeUQ5X7utB4MejxbfhB3ANkcAOYoVyQAQEQEfz3qMDPEgGYiYlHSLL
h8kQbEzp9zGWYN5C/SWPIg2O3CoYKSmtVzGw3DoyL2IsuuZJJXLakC+m680nO/YggJTfG40haOQb
uNqncP6Oy8/I0Pr4rGCcfklXaeQRfDNj1Ac8EmlDJY4Mgiqnj+jhqBam2ooTlibxLiBOTD1ZjKT4
5lsnMTTnRje+QeGGHKimMaeXztPsB58ej1hI7NC5bBNjALqEcW9GOhtvzIHaBazGpyEick9vgNhH
aZ4p9OlaWjDpB2zbLyyo0kClp6G2zn5oS2fhhpBrT9WYUCqh3w5tz9aPYpH6DK1J7L/FYUkTAxd8
fU8i6PrTFI66f616Il8syFm5PUAWOAULwiWYvr9HdkhkHwQUh9OH9Utgafcr0GUoZRk1YLSgKsXS
A/WMUnIzU3ux8MjiNQe4zQiUL3J2EymfND2GgOgFg95vsrG6ybBYzfGTcmbUQdq8E15RC8EWMezG
c+0gtmIR74SdIBVt9RDO9PckWnWlG0ZsnmA1OdrbNfJbG8fM4ATHF6D37GKrn7e3Vi5XtrSY3jD0
vwF8odgmKMuSXdGMFEJgdixf8uCjS/T7eiNXT3LIWQEbRHLXgaJqT+/VGD2ndZ/cm5H+EsgweKu0
U5WNlxdsKt4peghsJq5DnC/aSRVvuatD+Abk67hUUgGfJaC+UgOoKbYEzMAgLegU3A3GrdTNQc7O
/qWBy/BDec5tYtPc4wWvlsPjaZdA004ebvm1erUmuYM33P6w1rNC1Cgz0j3Xpc68fpMG2vMeDn11
hHhVPRc+awyv3vn980TUtKndf6+UbF9caxfMjlGbA3rPABSjBdAHV0Fp8QQu3Y82CYoaHAQ7HjVK
/vH2BQnHJVDMtGlQTpHgSjLEfIT66XWyg1VGdFgVTIYMi+OWP7yDAuSfDbjU+AdgVDUmpygdlOlj
c4mpiL2/4QKun0Fflg9uuCts3PrE6W8NmhpOHTzct80o2+DariqD0KDelSSmDvIBSzn4c8gFjMhq
Zf5ReCi0eIKcn+/RxrvPafXPJKsZR1aDyFJ7LudtvzmlUrCNWyJM8PHMLLsQc1vIcEC3HvYl/BT6
qTiEQfcDKirYdBX3QzElv6BURKDVw2H520YvKeTWkV+e88e4f5Bdjy9Reqvl6/01/9ZloZwucROt
iWRSF7Vfbv8rh/Z1dHOn2Mdc4UXSCePQ8AwKkrEkzzVk6qIi7w23Oak7ORy5Zc6aFw3gJN64RsZg
otW5BpkT8u4nzMYHtWq9DXppj4d+oEbTLYK2m5F5/4GnCRHeMr9luGwDCO1agMKp6loa01A8MCY8
3K/oz2xgdpPefHvrgkZfDeaNa8tKcyT34YfrL4T3SOzxa4rbdCN3PeAAk6dBpnS+Q3fzqMBjWFB4
aJpBxPPIBKojK/DkYem9ZIC2M+iCke3ds/+tmVnxlslZ0Byer5bYmLT4VKlR4Q59/xaV7o6G+O7K
bQza7jDsBGqccOtTHkZFBBrqnpN27T14BcYIGjBxTVf2QIZ8mhMVZS6MDs/UPKZR+qmQPQeeX+tj
vVpZ0dPzy5EiefqTZcaWrDKikKRHbfIwhZYkmVWB33ilVoUwi6ly7L7nYGthsSe67HNFgBx1xmHK
Ux+79K8uatlE989Gwb7X+OtXTBuo5XuILiKog5feF+C1E/ftczvSlo//pjQlxEbjXWU9UwZD8gtc
6CDYNi8BrcStl48agbn8THbm04/09oJVxFc18cVeZe02wIvLY+Zhq6AmmsK5mCsgJytJ05fpfQV5
RIYotr/ZeGlfc+3dELY9baaOH3rSCwnC4SYZEfp0Csuf5YrodWT1mngzLqOzyMfl1CP7J1eQbQse
c8DDP4RukXE+tTpwuNQWJEeKGAEwu9AjlGRe4t2mxNKUMtWxr6Mdg5yDn3oNYLz1bsGtjOoGv4it
SuUovGLKJOzkFGsasBjUCqC3Ex4YNVEx5M+FpPMeimhaWpdHYIUYPqV8swzrn6uCBD2UeeZdIZ4a
yxkooVXQMjo8lNAsDdTY4ZR8jDB2Hv14Y191NYKJAbNNIkM180K6u8xDJg1lmG+YsU9AGc5eY+3m
6fbaA7wbrtuM27bgbIqjIHe0qKfd/VqorvSOayYH4751gyYTNx3rxx8sdGik3ckvuZvvuiJx57FC
ffJYJlPkjdMlDC6jQeirhzil1+YQchn0T6/dDbJQAhSwEgJJIF1x0PDTvpijnOU0rW1Eenez2kG+
x+bTKbUCtn3lw3q+w+H5MqXVduGFpfrwZDJ1zNncT7BBTe1fvhDnpAReP+7buav+OO2WPUm9w2N7
oBqZnAI3T5bosDiq0i4tNAEk9W/LOcULfaDr4oAfRa8PZAG5d37ugmay4hRQyIiwI2wiDl6MiFg6
hrsUdijnqWUxocci2paj1smaRinruSmxRrynaZQ8/4vtlw3IRGObXYadPScvHlOnWbHaUeVQohAP
VB2Hw8Iv4XLw5hv84sf8bwJZp6vfxSbNfLRJKe87EltsV6lmgGh68JCuywOX6CFr51VgouI3kn3Z
DtgmoRpwl7tGZZABRWfKrbuyZzLe26zdj1EYsqSMZdP9GtRabbEkjlsXbKwTgV1CFs6kYNAGayF7
wtQrRB5PP7jwx07qpFTZKVYLF724qyBKCx/eCvuUt+e67xuRe4+IF7n8krhC8fgHIJkEtdeoD45V
OVDsNgswOTTncXJp6kSO4G/BY6dPHceQzgxcY/iLSpkdoPT6c5vxMOwFy56qsYdCaXI/HN3Bbm9Z
HWOgPqsJjRSyNszwYRabJsY3eCEGNCk8CmFeUEF6XxtbquEplcb5sx08YAgfguTAu44+B10u1ELm
hUuqxmQodscAwIaaZAuUkxMdFpWlRUW5c1xgiymP13H6HOk1EA/qnFJOQK8x6WZX4NUkuG6oJqsn
/Hgnff2v0Ob4o+j0YjGJGv+Z65gMtk8kJh7pASEZyMi9DmXN6CO78hfe+k+cOMpZUz2UQAKKGBMq
0RCrrM8IV481vaf4KWNV2IaD563z2+oT/kWYPnyU85PApYuOxlccB+Bd5qdq5X/li2IXD3Zc2YdT
MiTRCAY0ucKCsxVEbTE+TdgmTn0leCIhTMxqSgkJCNyarMrMCZX5b8bBAAuhPuaytoZ/jOFIXuPn
0TAc+NHcN+UtRWqyN/iMN7Ur7200eVoPorCae+nCRhtHpK8Cx5o4kqbH+eKfpxRmkKPsNzgFRjis
Vo+/GCm+dMK33/KiOxPBHqMPGrJBHRt7/qEHgoq+2QWxZtVWLTjbYrFtPSxX1KUptCR+dMqTOdJh
s3fn1W/SqvRi+sm0qHk/IKVgc2y1/Y7FoKOOK+FsC6VzKNQDwJ/x4seooUCDAjS7XiYSqvPOwqoX
XsjY9vs1fZrsaITXwcaBOOIEOY85iw2QqzgOg3KcCsITTpu6CqYLrVttuU14RpvbQ6iAWT3y4K10
CjAd+WsT9n2DIg96rf+h/kQb/EYhhaVr5ar1H7mIBUibKfLhvdKP9jp6sLD4eNUwNQ6DndrktaBi
q57hCFeiAjHMWb50zZmf4V7W36azFiywIWSXzqQtwnm36YuCUmIeG7qkyjg9SOnyoBEKnPIiN9U5
t0HlaVd1er6+29PedDFTKh7HJkzmPTud6Ml4215HlclseDVBZPf8D3jIEcd0BY/X+OnCdkrkCHkc
tLpUmS9JeJWxU9CxDGu2z2bPpBlqk+SQHPhknlVb1CTz/gt0z1tS8lLg3p9UspQMNdFca2uIf28a
N4mzxsn9iEsEuzURVS0tS+UgJWYouBgd3Bkto/uHN5me/eM+hspQnWvzROZnLEqVxm3rykE3wN1a
pqpLG+nB1lO3d89B3nExYxT9SDEwUlXqfTnSKDAgKJipeW4qr1gWkTVHQykt0YR+MOdURcH48/PF
S1V3VzG9wdsmsOAl0Z90/JPMy1+jmoMP5vre6DU21AKKToPOiRdbyE2dMfjjUAgnS0kZ7PtuGolz
J/Jg5Fki3G5bCEuyWEoi+8qrptDXiPV69Qvx8PRDCwwpaECVACVFWtXGwfslqe9rFsAzt5IN61+g
BOCVNpUeMCnnIIuUBn7+OfMHUhfZlJ4XohwVcAoubte7Rsa1aEsUwqVa5Ek8QX4c7FY80to2CI3G
Q8F4+pxOa+B4XA++ZYat3UZIJLlGlzs+wNuULzdoaSehx5eL3TS5ZseYeYwtl/zS+k/Dk/Uc/Ewn
8FG22Ia5zo6lVm4VfgKmD7YPA2MuQtQkrjTPNuSCbwMAtNl+3NVbq46Fej1q8X1OmDumIIF0Bixf
rWfLDndh+NMTxi3SkUTo0h/9Z0/0JVKD6sYNfqUUDxGIB5sHImXd3etTKZIDSbO5J2DRNMhXVnP6
V0pKljFm8x0j6Rfo3ODHc33vVb9dXsvg/LpLo6IHL6dA3hJSedaYFOMaCYN+iGP507HK8dffHwAE
dLINkGXlBNs/8JzZLVjahOpFqWz/EB6bvs23QreaMpyV+pM/ia1ruYCMDXi3qettbqd1BL0l6+MU
3pfWHIwPn3PR1ci+XCk+9BvOLaLqAwfeDKdCTTfp9j4mIvgfEgp8+UY5+TypWQ3o23K5zqMY/Csu
xFeS3zBUEcBjI7u0r3UR4vAhKBLCh1HnqgGwhFuXGcocSblOe1upHlwJk0NGVNpZ3cfziuRd9Mz+
IVOZeI9Cz1ZKj06hCIG9j7ACrPbRqrWhcnOEo1jWKJ24/QYHMh1od65Qs1Cs/RY5t7sKTiTrE3Di
7o6FH3MbZFuWFMotIfJ3/BaiTlMAjd2ps2hqnxU8BuFHIOFnCgQapjF6PgHal4jWBiF4oJzNAmLZ
lIJEjdx9Gq83IzGJ6O9rrwKab1dkwNhd8GzJquDUOoJv+Z/PR5Ajbwrh4sZfa7tJ8R6cwhYqQ3Aw
/4WgvmFJXfU+fiQnKXXUHwlsp4ftXQnOoUSk/QaQjB9r5gfdo9b2/9QSz3VUeGVRB0VVR7naeG2r
q8TpGg6imGANbLKgAnyywKFgppVe9Y17pEuBmHjZglu4stHM53I7GE+ZBehz77RVTmkKR8n6wB9E
J8L08QRUYYlYzdaZsG6K8f8H7tPa1fawoeaaQeuwdrJcNoGhikjjq57Rcy/yMri5zoHtDDNBP/OK
Xj4LadRNMvWnOtNLd13biTeuCvPPJ7iIgvnTXxFa6KsFkhIIxN6PKDBWAD4WM/xP+PvEvB4CQ/pm
A24czjH5zpq5EiVrhKl+oWm057cPyP68Cv1g3mDZUEbiI+lsOw6/IW5CRizFyYR4/M7Xx1Owr60f
QuvGPcPYRb47bdkv5c/0Iz/AGAazgFmlIJqUtF+ggAeQI2k+HD+SrY8RqNVg0xLc3PkkQxFmOTUL
fmMJubc806pbL01EgyhryvYV8YFZqUIHJRl60KuCmoSmYBg4JA53/b5w1KaXXW+gEfkC9Dh8/4no
WssqGozN+s7yb1krdBwD53aTd6wA6oxfnWiO2w2wolzX1XsdzW0opgRCeJl+WQcODok6fCpY0zoG
DH03uar0JI9tZNYQ+VbLhsqdpVzxrztaaVvE1a/I6OGWz2h8wxLSKH33M871ah14AoDahgSvJ6EN
xtbeAUlW8dBc9xkgIsCRjBw1BgQ0VjJGiH3IpNKxK55j8Cqp2/i7+Uz6qGc0kfzQqOEV79Q5yfGe
8tRjNsKKeqlufNeMsYbhbVBlYcZCu86rSv1UlHHJNNo4u3ONMtfD7ufgw+0dwhJ7avucLC5Yeukq
WSb0exSJ6nb6CqjhnYwKmsM1ump3wfFz7jqAZP0ETJtyrLj2ByTclCgwiPjlQYYmAthwS49W6xqh
EuBYrpOy2S6sD8VhyLsOOVdTKAGf24/R95YmIyb4R8uVsZGd2CnwdJflZS1qGlOwhhYC5/w+B7VA
oMlaNyf2keF+beJFcOg8/rwTGX784BMoO/fjNPD7/DNRk+tsUh40apozPcjKuprp3M+MEybMWQDk
mwKltbz0N9q5E6YyIb8UnmaKh4IzdbbOr5hFv7j1tctGww0F6cv9QyApLVnpXZlqUY1K1+ea4iI1
3hY3zOQIZwEZSHiV9TQRddXp9kJhOCKIAPMGJ8XJKWl0cWYcbtEY7zamijAYdCphrhTlDVFoSWJP
/dIH8UUBkB1wgJcII8/rTTvhPYK4pCJ/eE/q+5H5XlVxXb2Da+mIj5SsomCi5vrOyQvAxPNzn9Bn
VwEc7pNI1vDjZSiJvLOr42f6Ken64BeazHvXJpY4mi7Jhsf+T2mXluan8rPozV3ShSBZhNc+xfoP
SZnOuk0cEMEGVViTjPQw3oYikd1IQNjlAyzBDSDl1Wf9RK+PN66ziWU9uNwYGdIQ9v/hZUzVyuY2
VvI3odWeB3JrJQgzGUkMQ/8XsnY5TO6Mmmnu8i/pgaj3POHBr9f3WnBtfQpyDa+gTj5Ccj6rUoDe
xsnZh0gzCaRCAvQzoVHcxGEsgKtuAsyyqjrHJOYhNIVujZAz8ljAH++kRxaH0udjxfedwbZ5ateO
4KIyfjgehI6KGc6kLoPq6Q+GyGsoqyQ8SlY87gH4yl0Wu2qiFprllXeLI36qmSKprPOoorLgRDXP
+tyxWI0JUn1zdlQqZ2qgw2LJenV8D3FwSTzfe6kYK1gPk+FR12ulVsPO17tH7KK6qto0AJavkZ1I
61Dnwho7ylYiJ7+aLapBfiECVQLp6OhNQHKCGsgvQtM5g8OFUfw7xwwJoP++CL/vmZh1j86auus4
TRsp9oxeNx07JFnb0Ucqdg5Zzx2JvxqgWcx4dfNhsUr5EEHs53NMGK97CcKRDg/y24HMA47sp32/
1IkE2wWDla/5JPV9197iFHV4lxH2lYuxS2osqPbxd7P475AjqAAXAzIwLGH5fZ/R+147q5Wrzq/l
uAbmD/c/QOgOXwxI4yOjuLT2p2A3g+z5tmikjTLu4HkmYOUOtkFaPEw4BeQp4zY08kb8b1K31StM
Ynv9crfs+62inpKrItePBIUVH10dzE7HXdFXBe/cvwbfZ1v6acQz9UC0uWdxHTfkgmhyt/jFz8pD
QfBqhfqniU28OMJjFIFapZYL8WB9v2QN7R0tCCmuh4H+rlHoyQXz4NK6s8IliQChVu0nj3nA8mFq
sQO2qOD6sFEFz8zgXMKDYtK/XzHUtlt+a5GRFk1z+j0wJZWc4suZlezFrxcIqyNdQH+idV661pN6
kasfVhc1oCneU+bZeVPUE+6Nm5PjO43SBZnTAnU9zrOGkezCXt+++MK7xa/PK5QS6gb4KFaBw4S+
5mftmj4vn2QrDIvXNekWSxDbjCZmlH0l48vuvjM5fWZDTkDm3LatVSrQqgNLhwDcqzPsqrJuiTQv
wJRVaijqJbgNOWO93liwGqzux3X9sQlcvcy46V9/XfBYSv5GiOeSzZr6x/dfLj77iHRKEDbplPEY
5U9GzZUopBfEmQK8IIJIW8oDjsmddSC5wOMR7JpokOuY9tHq7TLojU0aO8hDktGmmgSxyQREKceq
5P9xLXB/Dhd6CZlIvV4n9BPQJv4gaVegSVoP8oUkvID/MNhzTuChhMUhEhUY9CIxIhIkE6r2ty7M
0Ec//qFwSRaP1NV9Aai4V3ocoyVepfnkjYCXhoNZ53pyK6BmvHAp4iVpOAkZp4kb69egpdND+ifi
3YRF9mEd4dG793Wdp9Xli6w6FqL0iDit7zV7ALODVnolARKkjofWde2tHJLxaHXj5TxRt63HJFEU
B/GwvuyLYCJKbJQb57TdWhZNuadMNdZaxZsf61UM2j/stbArRNIGiwMtefYfCor0pT2bdXSCmxCS
QxRh8Rhcqcvv75ZFDb0ZwcQN6018GCbRdfmSft3ewSbxMVBnk8atdLP0OrYRH6P3jjyWzEi3EnnI
L9E1IWaWYlHvZZ/xIcW2i0gXM9yKn875tMIPLe7dk1EjDsIIgCLJsOi68uvbLQTDlYs97m3SGPD+
LtpPvQ5pEJeX8/ZKIK0VLKU2KfNxZtnDBtb5CyLBh70z9n9I6uWCEh7CV/nDEghW3VAIFJE5Rv/i
lxIm+H/EAw9OWbbcvuf/WXQY2jlTUIzxPK+JaCl0Y2Ib5U838xD/bzKPSayW5hlTIYGDiexHGYvw
FpVlC/w+kC4c9UolSSFjCAI9qH6wIK0lmnF5Wd1z3zmB7md/oAgluF05Ya+Jc4l9yg6XGRBUB4YC
E0mJFBSBKPvoJMm5lFoXmlbk+7X3788Bq/IshjT9ZNS1kAARXK8um46gi4xysbvUK9CM+3H/B0RC
Wuf6si1vdEFeemO+XssREEcqf+HdmThE6oRUI9aEJo/ibUEJtsxZvlR+SpYifk0TezvhG/EwlTRQ
XddsL8nktzXu2B/h4YHirHmqrsYaC+RpwELw4G3wgwgRPoEtmbvdKwE1Qnk8014G89NB9lrrdsZS
a+2x5sIqXeded5s0W8bDeUwN5ghWgogVSaAxvgg5cEhgaaGq5yR29xmPSIhDI6INRxpuoSLbA+mX
4BXogqWpBTQLPjhVRSPrJBoFnDRqCjVS0tuQ/xvOh34T1BEd/avDz/udWYKkPrLeP9Fw6szS7cC3
BFxywQNglrBFR+/b3TFoglXZ/wn6pGAmbwNmMMlOCqvwIawaee63psNP1wWODobe0FzMtA7E7Ejz
xsBwxmx39M9A8+ZjWwboRPtCMgobkTl7Vwyw4yEk8VlIgptTwbIphft/nhFQ/zQWvXLgquuzF04V
jKEdOAgiarzc0EgISCW3fnPBiOa7GLWsXUXRKPkLSG90YE23iwp6HWKom039qkBoK6LdeoC6NJj/
8II+1/4YBLMR+H2WfCfNOi2W+iAHIaRRBlWYxccC8Xxjmv3irViCNbH4I3lvgCX6Idi1RFnrjS6M
U3ZK+AXXqtBo41qFM6GBWZOPbj4iLz+VGes/syF1VNmqk5D0DuLzC/rbNw03zJC9IIeEbtLwe9n3
HwyXFrwn/Qosc3vIv/lO9DD33kbqq3MEYe23xmgiYNHkTe7cckV2WVgSM1vIRhZThBquB1E4xftg
E4xAVY9GYfb0ceubztv2Am+RDg5teMgW44M9l8Qix1NzA/CY9n3Ddw0m+GJr/kmRaQOK42obauXV
gtS7jyOwznEL2pDSuGEzLTBNgaA4KyhwjtB3z2D6XzG7VNpUGeSfZirXtUTGj3aGsmT7VjxpPpZV
zESTFaOKxsBrN1rYuQNRXGTBGhGT6X/zRrcdEZUsVDNl7zVcpI+IY05xlA47G8QOJ5BmGtJ/IP7r
0snbHpD/fp1ACuUPmOIn9TLWmTBE76fQIFTdNY1VGwUDO2I9Lm0KsjxQuLZWDMwm1fu0vFwLPYvG
vp/uhvAUO46Gtco82oxMhNXYQq+y1j/fZRHreJTkxqLzIkxlc03/qcclAGec1bWTVmMWwer0DDRU
TzSwQGN3wENbKD4Gfqtk7+YeesETp9uJZUzOmr3R8g+LFJjLNiNUExgBSSDiFy7AgWwWTw9n7kzd
QnoQly8TJE6OUv2a1EEVNp6yW71Tx4eVjY1OtbhXXme2/644xdo2NvVt3JDp0Cs4+wN/dfvJLCad
+EoETZj4dPUWms6aTSoQGlCV/cQuOOLy2RM8O0r9TXxqvO9+hXPgDmxz20z1flVJvyjXIY2fFvBV
7vpNOm29mLAre5YqMqJG8t8aRAjVW0f24xc3Tx2jl97GsrJxKrcKZHMtNL7sfM/fQqkQlSRZRu4U
VND49hjtsOjZ9ZglF6SisXuj1Z5ofgEy+q+vsly+A0ruvfPBSFSo7F9mWmSaMz+s9Ll9cUPucGpZ
uzrm4R18p5cTxphRR8nKxnwR6fP+F659VyD+ZVZXPmHzAOjMa3ELAI3NdFjCm6QxPysI2maUrf6X
sAY6xfc6By/Il0Kj7tUt3JU6WCEpwyLpZx3pU+M5g8SpzgekmnH1bC1Rqg34ruOmJpouQI+fhiDJ
EOdfHc7ie5SVWlSVZGisR1axGdEHlGxB8IlhzQtnOhWX5tQuuT5zdrCxPMjtBa1Sp2u+UCqu9hAN
JOWCv9D+6fSaE5ETOikzzmQW1AXFuVcS+QUjFs0Wpvz/Wbz47pPpXeoweQdWrvtoimZf7yzDdhpI
R6lTsSIkCYGNC3TajlQnfL4mJTuf39Frl63dSbE2SM3GVkJBq5/pWR5oOfNxcDKGBHRiBYo3e25r
HSFArmgYpBcd2e0VxCtni3/Sm9DjSIjnwqUjY8RmQEc9BpLTbCZ84z4lfQhTAYFsJW8iBVjNr6X0
jDa9bJS1U59ph7Jub8FI3Yaa6l2U7dfbWXLkud0NlmZxWEIUFiFceUZ2kt1si7zqF2O+pUvqOpEQ
nJ/qtNTwusi22FVcBKuj4fKqucI7aFXu+i/EXGnnpkLCk+C/o0bB2VHV0BXiRpOrH4U7EDUmPCgP
Bwzne17vTUHdoPpydZg7csy5k1K2llIkRFLsJcXfumsl08ChMlv48iFScTYwlTv8xzulU7L5wj2X
A4gt+DrvVPyBVaYFzjwpJ/pbYjvQxKwVjWmexLOfCF1TO28GAIUeeFzyPt2cPXpOVlZNsIoo/MjM
YcxwC8GzBccYvm0vtSYv2y2bSHmry1xlRLL4Gjtcm7WJ/GnsOF8Kwo2a0SG/Zyvbua4k2vAyjhNT
HcKaYD2f0Bpn1tUJQH00FSPInEk/RnX+03axSpcbIDmNIk6H8eRXoiOw0UN41RpOm/ktjM9hCwfK
ejt15TYSZ0BeEa8xLZcgJUDmZ0b/YHLY/hcyejDQGbI9Paf9XYGonHhC2O1CMGJN3h03BcgouyzQ
BoLYPkMvInwuwGS+Qn0HbfrViaHULogspMpCWsQBHQmZVEjw9E1bLPUl9rrcPl8NFWlzg4fIJdka
AXeWgwMs15cAeCi503FJ+jM8b43L+I8m4Kw1N9j7RzQ0nvBrx/K/pofuga7Kt98wcMYRBJ/lDX4h
2A67jIT0WTQyAtFKupb+pG4tnMb2V0FERnKyUQA7Tq0JLGR7kwmekdkI2HLGxyEIHqjKAUuZZWa8
vOueikfnOGiYQ2/GTat8QYqWKzqEO7Mmm4Y1AnLlvjovev550eWcSDG3aJ6g/506kHcvZVhFHWnD
aT06GPY0ZNRgiD8a9ETfTzSgPn9GWIOVUwn9gbwAlXYfXJvlo900d1HkSuSB6M+WYk261EY/NFsN
SK7dYJd1ps1nhRajN1NhCESS/ylRk9ZY/lAsz9onmyjHSzmRt5FeEknrphxshUQUDKSQ9z1lwCLt
IlcFgJgMlWqMqvvb42IKlOP6HvXUdvp3LLqTqvrQikXRsm8m7m/zQXd9iI+de+zHu3R7rBNQFPns
EpgndwQwZ4gNgN6DPiTB+1R15A4p+U+atVSOqftQ8E0pn7korWu514J8fFGUSyUNEm5LHomDrJ3X
Qm+1ApwNq5U0iR1/0G0J+/oJVlhLBsBfeD90iz6lSqzByK8hAW6jpJTtTaOyIDsijgIPpqY0OHuH
nvruzC7XQX9F/rMCzfBW6KgzRK3fxKtfKp6RmVZiBNySYn/h2qtmdbnYC6nXy2EGv/6ctvITXCCK
R+c+5mokB6O3wJC36NP8tlVHqJ4LPPRzhXGL3ckfWTW7cN0QMfP4vjZ4pzEG5Y9OkrRqRe0u3lH0
f9VirfXHLG3T7iMO5MI1biDX3Fs4pSH6b8BQZB0Rm5wEgYPqOMJBTjkjBlBGaPOPus+w4kO4Im2H
hD2BBHxoXT+jBAt7sRiQ5fWQzCL8W24u2j/kM/9p43SLNRXyyXskX2NM8nuOvnLs4K72uy43C6GF
ZFdxJXMaiDR9HKg7X2O77hr6NFJ48Iq6d2w9FYiCOtw+qHcdbLr2Vet+UBRxNObUHKDLpcORvw7F
h15pXOf4DsszU/mFh9nq5MxBjsa6WDIS4EcRqSrU3x21niui6O2QkbE8+HWG+OquisS1IGJ9XSpx
OztgGsgzI413hG6jMqiWKc7L/1NDcObCyS7R5q2cATnTFkmhNKKDIJt1PkFt11YT7qDk3ZL2X6uL
PC71HHVVyLviQuh4OEFFzZDWLTObVN/Zevu0M1R2lS5oiNgZXB3kkVumaX8gQadj9SekkPdrmOq0
phTZRm+yOPnvUCBmFRPh9g29iZgKQzB9BrVh2Wsbj8RfRXNUVLeRnX8PVsw48/HwdRdiotrx2N28
18fgUN3JxA/Hn9F0vLvKjDPnMKc706jr4UtVHxzAxLcoW/jGpaHyXjQh7Xd0LosLObjaIG1rrlgV
0iZ1+x/cXsTVsxfjsWMYlYU1OR4Nybb0VDKY310eVpsJlXQ4qM32dImsa8x6IDbNKisGMMR9x/BM
Q5EP+JuIip31mC4YDjaOHjthw2Ayr7B3eRf2dAmDbFah2OHctcpaAsiaMANSaHSCixxXMx/ZL2PJ
JOk3PMTOZyw8ACGaCzbNXVq8jN9nM8U+DpfnxwqO7ffXTsZTTGgahvLv6MDZ5NG6j6pM8iqVMOkr
IrDQ4p6adtbsMki+35Gv3AaBXe2IBYYUqEIn/d1FnnMww68LNxD0+HoiPyKfnlKMF0R1719oij0V
kLk4FkTQ3yQzDNPsmXcqq2H+OeW/IOPEqyjN9wHj8ZlenAkqumfHrRw26L7hd+KzsU7FmgwAAqSy
PEnHmdEUyQs2v3p/YcMYtyt0cDUxX6P2PyUMsN3ZQUGT8ij6BqU1LGenL5oKqUBWA8tdr6K0ymqH
MN0A3/8d973ISQ9bSGS0y2H5Tx2a5e8PeXqTrzEkqAjcJbV6JANj0RCXJKoNHDmlPR4XkHlQqOVd
XYlq94IVmcPdKXU1qGHHUkzUzVdNoXxMOkzqWljur8/dv4ENwz4mq3yveZZZjdOYzX0gMdXkgwGv
NgKP8xLe0deTsRIn/6pmhcK8gYoHWIGUYxRlD3hAsu5Se2rzQPvhqMy1D2shkkmSdvP6gqP0LQQh
wpTjZ3BGF2epBr8BRfdZUxCGyiXS35iuwef40nA+R2/UsBDq/sD+NFaamtp+kYpk+KC7Jz1y/Ail
oZr5bph6sgyWd1t89u/K2EZZddrhTKB3M9gpVY0WWcNXBfZxDgZfwczhB2hz4cmfgQaIXvJf/5yx
ZHMhpodRxUDujaxJBFIaGaZvr7Yu40LSOUVbqI1bNQdqhw00AAlYp9OXFb48robeHJ9ZudkbmKwC
nmE8MXsUvB4TRQAW7UHxdIhJ0x8mgi/ntdDrTAnOBU47A1BGQVS/VBzm4W6eleoj/aNn4/OFv8m/
zFxxG+/4tzcvFBhLKOEIc2lZ9Ti8OQIiHbOMDzndEWstMLnzniKc+GXMfY63xIlqBWIM3GDiwIT0
EBUwDgPRrK0PEekZwYBL17Uxto5Ayc0f2WM/vUAEzl7sssCe5KSTTF/kdBTL8ppKXAk9sCwauSSf
p1JwPoP/bzOCCIA2Wr8FxZxD9JIZUTRJxOgD06cCzoe4M+Z64fEksSdz3y9oYKDguUHXSle1hTF7
hgO/YVOB42HOQa/jafF/p9D6ZeG3S+yK45QuX/+SyyBrZDa63gaWI2fIYdWWrB2sU71rHcs8Zar9
+YmHkRYnEiP7sQ0Kw/I+iKL8GJBsZNzc4/GcbLSP+/20wd3rV/1dS+ih/25RY5gS9m9ywl//vZKz
CHVFFqbqyctmObuU+BZB0V+Ug5a22B4JBn2L6SC8rRJyWKTyykiBi7PHHPOkMoFidPyD0peX4bNY
LiLULO+JKgR2Q71+B3GgHxCIUlPpzALRbKP5UQAuc0l43ffNyR1Pad8F2ogodaILGhxL+clKBANs
4w+RxGOFFBB7s7Wwt88+ZPrtFDl1REK4UVrsaCDooEhMjS54ZLsaLL1fJnDnH+e1JxNdmYnBSxLz
OlK1bSQ7ecGSpBm3hELFE+EA5LMS66twzKUlp+20CS1LanSAdxboC8Y/ly+ooqeuodnetBeVBmzs
PNsDtSZhU08fAIaK0voC2U1T+KbqfF85ja54BD8ad3/sP0k+mJnGf94fk1SzbHF8r7ePXMJjdU3c
DEjuvshctCrvqN+FHEe/t8DDVg5BB688RG5knDAqr3L4JuNLSp5MVK/Zjp+TyNq38PA/aQ87sh6L
MW3hy2pOUPTbq9Vf60hiUgD41A39r2gCwllZ2lYSSReKAdmDV1krfYqI2xis3ITtQg9qM6XqP5i4
q/BuDrFlxS10GH9u8kyfZYq7yQ5O7f1AcoUHf0+SPzApc635ccDc9HhY/76lVypZ2/6vFz5VBkN4
zX6Vf8KZof8Wk/k9JaUzF8nPR2hNzIkQwQVxtisrTLT4GGBpVbkunN6QzuEQsuJy89bKtjSU2QTX
ENU5vLBMXknAxhLtomyEtgsZiyYKGNHcyGnSyXnZ4L+5ZFH4YvJ0YBnrTdmcAQsIXzB87DnL76nv
9k9r4WVq6YxcThpFSPFTHv2g74DhcWJ/xAryisHq6dnYx6ItO2K0KVVbqXoSR3paWAkkukIlOEHS
gVuwqGb02DpbL6roCoE/Za/YNMsiyO1K0sjDnjPt6v8R2mB2QuqNJh1LztPSoTnpjQpK234FOPgN
8k9lVUORADnmh/VjaKUt4mNAYwRdEK919aKJZ1roVOv3+HgT7KgTOB04VFtN9Iiui6ycF0n1dfYn
nJQSm+yjme5XkmBx+4HQC15VDGYaDZuGuM9mUY/J1+iTxsSO/c6aTfFgGG4yX+4sxCpdd48hWK/M
xnQmnF+A696yVlLULjMZmgQMd3tIPrOBsvAmraC5XykBBU1MB58WXZo8d3IZPU0JdoGnFq5ipIoW
N1SYd6z2+kBMk63yYjHw9QWL3JXKLOdFsjiVXRisKzzNW61V/wk9q5CNzAoHijmcUBdhsa0Z0xgV
+2f5lzHA0+MCV3g0bYH1olZI831e+ZkzDu/qMU6eCmNn+Ye3MZZx3avoNd5U6oqR3lKw8iAjkMzs
JdAAUWOiVhKjowDiyBn61iO/boQmmCueq5XDs22YdtNr9pMG93rcWMDWSCAdP4T6mHBQiCeamC3D
8fuEUXjOJLepH1I24r7ofH5yiaujOheRRvXfhOqP6xas6gb4DtuIUy7dZJGVjA1rlVXwJ4sa6vzF
xHcNXflfHDN03dsKqPOa7K+27nvziv/qHJCY8kZBHfoTyOoAJv1fHS93+L2AmUUIvsYa1RqgM46O
YHBrIoph+kH3cI9mE5vz6vGlFUT8HEDUW36167bisjg/DcJFO9U2mH8OgMTBh7YJbxVyDgAyi1Tg
4n/Ixjt+DN1ImDUDkD7xgUjWMWEgrEmrts/jFrcgEYC1Dw0iU6KyaGrUWpsrV1XQXe5B8EL6DhDH
imjrwGq/5uPdzDsU1Cr5ON9tur2gV3XZU8SWGAtiUr1VJKNC6AplB4vQZXHcP+9GfLwep0/3B6SZ
0yF0ni4WeTkDvrneFWfsIBvXoWQ93d+UUHo94kBN9JWB9pXnMUbuBsdQ7HtKFfGoUJeN0HFNT9sE
D38TP2aWnedynmXO07RANfp+Da2KMAmH/LYmxwahHEiqy58cvY0T4xFrnfXWBzksbl9VKCygaPx1
LHE3eCrZt/zs+/96BDKVgj1YNgpvZAEBacTPI1eEyF9i3N4+vddqWQB449wDGQrDzsOEVGM4F2AV
ekB3R1qZ9q8ZWaHl6Z9pDTyS+5JRAKzxOW0SFh+5Hns8XBIhUKdiqoqds+1vu/7XCeIiWHdAp8AO
4jNn4a9V6ZDqwxFgk+4NQ+1IoaLlbVkzLthSu2z5mxn91X4D8arZrlSDJya5qDBzMQ5mVivylF9+
GOcXnKtMKOswOklGzmIVm0imSSlvAlBcysa1win1xv9fxeTUmMT7Gq1psX3tKXe6CfIQigxT6fFk
+1gKLYXoA6mKav6KgVPmJVFmDOhbJbg36DPjLgQcUoW1jbQkeYd3Vs6PXBjDoE2PrH3G9RWC2qNW
Kwzy10l91VDGzhQnpK2d2ozo7retVcqL0HiyDxzeFH4BTw4Swa38RdWHoJ9KtwWthBOfrV0jmuKU
+r9fzTn4IbSrmkF8NhpIoiZshmM4Y+ip2BBcODPzqR1DeQ52jrExuTHXGIyQTZmeGcv5foZc5oA6
3+C6AFukGSt8zGvBACqo7HJ1UuzlVmlh3OWkJvvJ1wnS88Lbd3wnQTKu5OEs3zfrCrQLcdn2sXB/
kqMq7ls2BGdlVDXakVhnxlIplJ2UaRn2mPO4rB8HkvIHr5KFBxJzsvfDh4gQkfNs3OD0uBUe8Hs8
WZyUIO6H35Dg6JrVsQDKb0eMDUT8MxyxVjfcbQLJSOvd6jSmG3yS0du/LKJrE1sWDzp34QDZAsBZ
GrwTZA2FwisiRYJgeYYJlXmMy9I3hN1P4nwJXISz9OU43W5yHu50cuouJ1MzYfqwjgT1+u9meaEs
eVIb/fuVLYz3VOQv6io9G6AECvxERVszpY1jWg00q7Z1SfxzHmAPfhxJ0BSPgB2AqNLLlOqdC223
Yw2fyd0zhlq0q//JIxFDL+xy8Qfqg5RoI8nanByXdGYsOuxArpdZHHkKMwBbNbwHZQq5pNU8a79K
FEvzh0X8CmrS2yK0VLVRX3YzHRNaM6wNvAIVbtOth5X6JRH6IWb2akKmJQzVqyKAbP+vmOrMw5GE
ACYEBl6TC7TWiDNbmLyIzlx79wlXBwzZdxRkjaMBGsn14yh9269wHKgBrO5WQpRYd/etboISEBZN
5yatB9Paht1SwzOjPlaqZdN5zRArtvSRhfWEf69T558YNOj0nXsa1ulIPa72/hHX7eEEkyI3qwsl
PQiYkNWdZEF8ZoeIb1eS1EHWTCD2XdKG1G2z0lw2WIqPMa6VnjWTQ+NwTPW9ySaAQX8WxC55JF2f
9zyifKF/OgQP/mGwzS+qsoSWlGQ4R47L8Dsr+ZOSO/LKZ3jANmwBcZFPcgQ3MUFz/y2qi8uu+Deq
umixyDTBj7Nvrf0wDQUQyE1z5nRIjxl61yJOPQXCmeW3gWAdU9B/xDQtJoKWvKTAkNaK2DjVlnzT
3Sjnwf7OOxiaklHVRzqaljrwzJG8MPnAg4i3wGxHdWoV6nytTz4nnldVqEPrEXMFTi2BCmLSsLTh
RtcnVAzzCjHDXUatLGkTuj9mFPO898v8W6BpNsrVG7hcuAenqrY+D+/vAZvyJTM1IJPOsQpf2iMq
/ZsaRWcrbJyjvgGHB1ELYyhv3OoDDKdWViXa7DQ/6I1gZW06dIRfjKTF2A/VsQ6mocduZ0GUAxc0
oQT6WX2mlBupNcwwKfnDpKWaeW87V41lOo4r9XZBXadxENghs2pMG1QP54MpDY9iHSSgK26XHxC/
Lc88+C2SoIE7GQS2nd+xUjyiYgUuUq5zp4Akve6Qyeg50P0spNhajiDd8Yoext727zyPY2zifEOl
93Y5yqtnG+ImJYGPSPZc6eJaG7kzJ1qX1MJHiNPl8YQzbDY0mRkRFOUSd9nzoKDDj5KXYOaSKKL7
HjGbjoAHTUiz0Tj3q10oKIZXU8ZU2TdMRH89hLTjvfTChqGASTbJnc8PxsL5HFbVHJc/urA3S0AF
p+YLMcBOcKtTJTaAdFVCjxHDZ54qsYXuobS/YO4+hyit3ZJo/1NDYD0hLsyTnkrzlOt3QZPMUZpc
U5M6sWDKP6g8fkDuTi301trAAUAH94DBdm+JiwEgDykw8Thxx44sucYlRP9MDHSDaqdPunCb5KHL
AOkN9V/C5IecvERmbvS10Ruh9IsojQKY8DL4i4IgVfTr2PPxxOhgLbDNKrJqcQBN7tN0QXA4iir2
Z0RAcd0gEinzfNNvfmMaIW2wOgnJwWXqJtKtJcnTSiy+trWE/Jx263XVuhb7uYiKHvgRhCuC1jqg
c13QxIVV+GjqAfkB7NF9/4p31hjQVbXJh4D8lvNTx1Ov7olF1paDcgu/xS/w3PbvCPtSoCXldIjI
28QNxqMSqPr2S/QsI/33aydPasXTNygEQhibysXjtbYYeHUqPGxldallrsf+VCeQlVqQh0wgOa8f
4ARPRWqwzrKav7ENwGq2ZXp3lgUBhh4+Y6i9S75t78AzWciVegw9Ilj5bVCwlwl4qvP/8WBfPGGf
qD6nhfET7EIcR+uri9TcNT0+aCy9FM/st6dJKdHWFH9MQzxQpTd4lhxO7Gr73wmQmLcgLggjq4yr
0KNOAktdH5Vtp8vwTnIzIZKBuN2+hv4gcjUoK6rQF6vk6jJKP+OVd4PvpCHu7ullJz7zTpRSgOn2
OrPcqX07E1pAqAVHferVq3zLe38shA3msP20Wa67dC9Dpa/JLgsbCaoClvPw54qoRGgo6DNw2cM0
l6LKYdboPlRnIPmnlqJiJYkr37Dgkvk8St2J3LGX0/ZT/q5A5Qs/OsE2DiMRZl/2vIvvPnemxtRh
yHrYr9fZnV3GDgI9TkuQga5m7Dzu7IMAtk2frnCObLwl8Xcz0+CCcEW0amykT5Cfij47XEA9odHu
4ThfrUfKcUJ4zzYHAuALQUfiWH5AjOStrCfq4uhqQ8HW40QRDkmbXWbYquAUdsApxGB6uYrucMmt
PlnlIvCQjC59TmGWbfpDNLUpprD0QnqtOl4u3OU6F34pBpUgmBRMpRCvK6nU/SICJ35Jh9J/HEbS
nNCvYCez/l4HACQI3gauoJiJieMA4nMkkKmnSVkYPifFtCKuXQTLqyBoEhuVxbJNqnzI16pGgDBS
RKcF3s0oJ3yCHJWD00E7qwJSwBg1o36Hg5t2LQpSOU3csQuqxWP8lsGD2yMuoaTBOiqg3iv/p7Tq
FHgf+suiz5MTVDo7l8uCwwpIYuxx/Cnv2AwtVMx6ZdK5JqHWWnbdyL5xIEJSzpcHWJ9kDp5/2mdc
HPCM8NWGzxfz3NjNRGD3ugIUTxKRCgF2QiJRdFBp1BKCnT701B4920zgIz5ueCeziLfVxa2O6wsz
5eI1MMADZEyN5+w8Q5ymFbPuO6+L+C+9VjU5ub0HeIJ8mvgvS+Ya1np7bjrCfZgKa4VTY5/z11d4
C2hxX5lHtAU8Nu7sS8Ez+gSPK0GRRDAzMzbVATzceO2AqW9dq/T9EKdoEoU6mnLjo6QM4LpqOmdh
U42pnVpn2TBmBUuscSckAr4frVuzpbLpywMNT44l3k9p1eOPsWRG0IiBkmKoPYVMR0UmaG4nEwTj
HhdYZKwsDRPRogQlfazZXo++iQxxnDLVErnlGB53XRUOd8ySKHSrIj0w/jhH4DH7V5QDl4bR7RYp
rHnNY4uo7c27XdgWiW5yqsODTh7hVQO/PCNVvHFbfLjz0QSU5VTPQ24Y6OnEsge52CQhWyH8u5MN
ariGnTO3+PqKFQBq55rmTg1NzRDLac9iT6YZ5ZPu+pv6WL+3G8KkGpE9JgT5RyuuZPGY3KAz2uoD
hv2XebazLlXNMNPvDgBtNGvdUF6tq/7guPRbCvVZr1r+eOZwBn6gkuXeYYYrZJOk2kBmeAfGXJL4
XD3Yx2mu8LT97RuuOzCx6JsmFgQblaZA71FIMVutzy6GFsvUcZ2fkXsAtvhAO6OKdLx39y4YRwro
wQaFVg3t/QrLjBm80Q3sqUqA34pK66ChmhdbsN0KWlFMsZSAc8wMWfEJaWT9+UIL7RKK+e/pPBYP
n8bSTwhe0mw+Rw2HIUo6U9MkvOU3xDHcte9KWxZSAuQakj0F4QSi/S9XvphRxEmXAE8s3tb+yWLG
oFHX0xAB2pcHFXCSWWpj5pljnWUYFvJhbNxjD41Mb4px2L/7eXzV0oOXPcPsCACn0RXrfoUQe9gz
3k+vrsE8l0p4mvFXFo9Vfg+0IbTcQMnznCPldF/MY5r8yCWuv/WkQCvRzVDRZFokNJ8exskP9shY
Enbk6cxBT3kFC5mlPF8dpvn18u3sVhznC1sG5JPPbDoU/85S1V1yTOQ2eX3AVbFeVS8IdcFmIXo5
hll7YaW5VkkfZPfEBjZ1/30k0WYZfg0hOagu1hS/GwlPVxb45DVgNKN5NwS7T65VoTA+Xknr+DwH
pftcUM52kZxtdyfY53HPKYIJoEqFv4IA0GDMVUZbMvEoZZx694OI1+SRLa6n4rKIYmlCI/8yDU0e
ov6emwNxh/yH0uTa9PXiZ4DO0hPsoVt5b+y2fPuYczURy5KpgaowRNjKuaf/plQdmyPqXR/XPkno
iHmX/eTJ6FkgaNQNNW4j3OGo4pxj4KxZtBgMULH1FP8om75N8LE+9gGpqgvcaoBKkzqDP+lByWDX
dBM++JeJsmBlQIiR7pB1/Z5RmjCc4i3XrsXjEEUuT9gKTt9MidMv0J7TtAx3QXI9/cwLUnss/Vzr
/XYe5VBL4tXuYlaQ+DBpfueFVgAUW6E2kZntW6RYnhcHqztLMLgCYfgenvB30DMuMtV5pLXMD3DQ
OzKKBXaXGPdqo+PII/Je8vmuUFA1cbAYtJUsaOY7/r/3p1HtE27tXa3VaUp4NSWsPRBgUclI4m1I
eiTUnXkbjduO9VO0WLcgv8PeyiQfaYHQy+fxP0GHXD6hyTjF0lTcLGtoHD25MUpX1OOwrJ7W+EhU
Mhew9wYus73pWoaRTbU4XMJgFElRGqxPEu/GTUQi2f/611DIxrgoLksDqQ6ks8vGpwmn59Bl249U
Sn4AwwE52HehOHsru4+DHnxVDrbFRdJBIkMb+u83zxFH1QeuoMGeupPU+Wcg2w8Ik+SCKrr/NWw7
XJ76LncsqH1i/8W0/mkY7E11yQM2dXv40ZNzpK4Qkr3AQxybbptaA5BuxTpilidRDBqtmLzgoiQs
jsRTAwHMqdVZvbq18UC4RUuSmlWyKD5SDftsZNQMBb6T17f0+hBV0FiuTEWE9KpqUVV8nvNFzl+X
ys1BIlDwGCp4k+64zPRpwP+wdygtvre0yp8D80YsSRs3jszMXtFdQ5Cx3Sl6wuJueOsJXprh0aWV
bUc36pAVsy5rhoXHFQy9764tetF+p48KUdwIAj/wvo+VPt34rBCiEtV+XOGCWpmuMZYZEwZwzYa0
9cGomABcNYxzcFt4pgYnSGtMCrFFftlpM++5egCon84Hxj36PXd/Lopsfg5A01OOy6fe8AmGvNIl
puFIcbJC1qa8C4cdRhj11Bjy2PtGwYFzGMig1ALmml/ftZN5GiyxEJZlQScxrZqUYO5l4YbWXXJ7
e/XNsDXbwwE3KWwb3DuJXZgsMXwAiCysDnLFaCme6bNbsxZqgsriPy8/Bf8axHwDPR+8ZU1+RpxL
rxdLzbp89YL6xxd2g0xoINqPA5O1v6Uf3uRP/TiU8ONJtkJ6yN+ZOKRfXlrEKSY7zZxjTc83cmdT
Q1PyEfO9H3Nf4MNH46ljrJSV+i6rLxrjR4mjWK5YM2Brvxe9uShr4yP+5sF/crb/reJb/rnPIO37
y9DREBR4RbUaxiWFUQeLE6puyp88YWRLa0fW6SKF2mQWnRHwLUumLtAs5zsfeX9pJ55Sr41czDJa
IkIaGhSzuTH937/89lQRMVeajqH2jKJD2xACGzg9zdqX1fXlZhEKV9FqCkJZFYV8LS2EB9K1bd6r
3ljHVj0PAxUNDN+2a4Kg9SOWvP4uolIVT00v6uZvHb0VQsJUbGQZBejsqmcqlE2DCU/Tdsk6rbL2
hHZ2wxs+uh5GEaIw3E1o9uKjtCS1eK7Sk9cZOLOdFBbq0db6bw7J4C3dm3AytKmoUDpiMafZpQUH
Kt1uPRnQQMG6yItRKyVr5yunDwbU8uCb2eket5+P6zUDLkv2/NriY8T6HMLkxb4WDVcLKYGize+z
VaasNe92SQBuwkRpV+H60X605CtKa83jZ90NKhXwq25AdUiQARNrJqqd6XP4OcmGctWbi0hsLoxH
IEIS4HAQzlwwAroZqINZdL1wjd29t/qnECWAhO9t4KaUU77Enmg5fPfzdyTGA3yxoW8wnmEZ4dn1
QbgaHnOwdz0MAeIWMkX7AFp+8x3vG2IuMQkoI+1ALeeOITOjKnJ87JV3AUCR683VV5FtnxInehMt
X19tDmGh5Bm5ac1dt/P3pSzXCwFbbn8ApUrRfassNhxwqC/+4xeAgYkja3StivcQyoyXHa62O4mq
PnGBFJGKVQqxN5+8cNTB/puc3oBCJ7yYJ6gjhaYo1zpCRgH70EgYmkqQolxZryKVY75LB2S6jDDY
+L/P2hy+67czmcIUCQqGpoF20hRuZrbAZPgboH4wi8ze6hI1pjgsXZyJSWUMXDmpCl1g/csrROpu
i0YuVPCEZ7qreabwVVNTRzUmeg3VRd4CUqzHStEJS8EcmBDAOfkjBnSyDc+1Fu3WEhv5nL6sYQcw
YQ0tGyweJ76YeXAoNz76nz/MffD4JHYunC/u1Vibb0ZrX19s+PAETMBlpjZqnu/NBtUkD9SWdqO1
E2xoKgvTlBwUQPRr41fjPlW1FOWa9f3sIndPvxmi+wM/Q+SozLevjdIbJXbYJb5UwQ6ynyMEJSPR
YEcqTmrVsq8jf/1s8rTXQ4YnE56OKM2ujkyuWz5DR75GPdZJrFBj9uXGBb3jlH3JZFXiJFH8hcGa
xupNeXPQbx7ZPk5X02b5IYXMQ4nuo36XtKe7CQ/EcsGO//hVQdA2WkCeeUkFiAVxPz3MPmvBGAUG
LL8sLVUooMdWzKPMRpFG+mYtlnam+ctT8yDRRnf2BXYtuTdV3Oe55yzv3k4IamqUvZfgV4DyhN1h
4NKjOjp/YTQ5GkXIbS6EUsvj7yrcHNq45XMZUPf0qQJ9NRX3bI/CMEgmdnCrrgiHQ9Y0n3mGtFa8
KTXiNXH8T60DmLekhAG2VVR5e2lXVZn3bWQhkwtJ0g0wDFUrjdgMOeTKJ8XbL/vAYf5SFuCGKJc8
me3XeWZbGdtcjvEwkk1SXVHJNjTUbYWA1zNHFa8ltoEUsuiBVy2/sIuJ/2wNSJqrl04WdEpxukgL
M+o6YxG4n6bf43906W/0v+oMtbTNTpFot7SXHM9S27kB7kjh1a6vkIPcAPVckJ0uP1V9uupZdUub
eL3j69oVAw+zSq5k2kmZGUDjZLlDATVyjQ5tOBqlNlwQEZKff2in+2d+6HdgCpTHrhHwHwKkknVJ
OAxrBLQ1s/YH2BXglQSYsWJ6Kus4yNEVWMKBij4Rq8O6xXrg+M1txQqVCAnGIBvA58iv+slJ2+mD
0O87+qOJ69fsJpOC6tcVdUaGxbZOQ9ldIOHqeOBt7QDbpgdAnoAmo0eV7XyoRWFb37m01wfmmZxu
E7SxqrW7nrFWHyj+XAHHB3DbL566Abnp7YBYkhaRO1iKX4r2om1suPqobDZy5eOPlVLPMeiaZzVp
4wLsi0a0rL1ccR13MTNlFGftsnx5NIRM9Mry30yEeS8sLxAusic8oinkafnFSEf99Byg0z0XTCKe
ysDTD8ERV4pSJrnTFZbWTHeCWFTzGTQy+XpsRqgpkRlkWRLCdewK1TDyzyOSz7smeFT31NrZV7Dw
kd/LRurQd1hVQR/34NMaNiydnm7Ck5Br058VuR6b5D5z31vSJWG3wnYCKzTYiqioLtMlcWcn+3ks
/w0XxvUJ5ulDAIDkK48fC4Gag6LZ/IHW9U6PkiSWgelFerP9ulRhMqA/u0ND2PTPGmiUwJJMqI3o
mjKEDnI1YB8ZpyI6U5Esw20ouCNG99dAz/GAm0H4hUck2FFj7MfVavMXCfY8Sr5iy3t2ESL41xAF
REb/OFUp5Ci9dhXHtXEoEPxGCNu1xcUzscMvwuxXr75nnRVWf90Pij4AgONIyXN8YQQx99tk08FX
s2MZx7W9w9JIxBgLh28beyJ/P75Qi5LqoOGplcGfR1+XEB459cXff+k0u+FbTUHsb4+omR1UYZTW
yopspJj5xcTx9db9THJ74yp0x+YnGNR7Jw9rpevqr7Wl6DvDtNQNY2HzpsWutVFia1xbQpRB+PW/
ZpJdA8P4+IOnKd3brA3fNdVrp38FZwe0HuCHdnMR+YYxrOkBqtqvlJfwFIQtXuqZjzn77m6JoHzu
N/FdeGftyg2rHN0dNjxidp4DUjGRmp4PJGOg15/CPPW/vrIlAfdwp2AmatEXz+DyYx4zFkmGJm88
uv43RIjxptBUOI3gnWSuVen1Na8g0y/5vQ9pXXnadABQOwPEby2UuLVYuzGYpakFNXd6Ed1gSvX+
+jcKzAgVHcV/FVEIV9cbnV7tBtJMxKiQtzCZpNzlG6quIC/kRu4ZV5Z7mN7/aNJZMjqBfVvSwrUc
OD9IL7cY3YEVDm2V8fXJFqT6CoJ1MRmLFszvr0X0Q+MNY6zQcKIhSteKZquyQ1R9KXyrWJJBCqHx
vQs1hZg8jQiEbve1UNBwu4rJVlYXqClGuyXe1QrvMUzFYylDLe5lNKU+FRHA8PrhJ7Pkn1uk1U44
ZCBNW/PD37EfMEmUpa0p1hLQVnV/PTCZEVCjTSDA3wQS6sO1Y2DEtqPyJvDkV1dApo2mowXHlAn2
XsTRzhGsq3z9PFJC0ZgMccmstmEwcNLSsG+DrZHM2DYRO8+qxVj0DYRieq7QgJUmjN+diYy8wUln
VyAk4iDgufyuenweLUP4hna+osy1StUrShbNUl9D25U313IvdjtRBrzb+vtNZSgrEBPso3gApk/m
ZOxFA1mVPvBjMAxN/KutQeE4QhvZQruKqSWeLA+Eh/jIQKv2RYGzCM4ugOL6DFqSPM9HzwBOvdAP
FNEa6tik548fnL7dqciQGDqa0WDjOJ3SH8NdasixJm6AOeBTdjJpEywS52j4hKmRKHVe43i+dWG4
X4T8IqHRYPrcsUARJn3aLjSLhnwnmwbIrdrz6dqnuHH4asAvrJyZjPOx45LEycxXL9nbs/HK1O8k
lNH7fP9tm9lnt3EszX0YMetocqCk9VQxiFcY3VmOk5FwR8zyLy7+DxB1cbkRK83VMkDHrUI3oajE
JOhyq3S/Oq3olkUr8eaIl2HeT4a3Po4oqyw+D0fWe9ydV2wjfycvgWXuMmatNVxKN4N4WQKRJlKe
8CGRDNFhkQA+qWxzJlsE3q679AOgwSTWTljkIYem+wpxEySOf1udprbx3BHFtCqfitPqmQx4ZGrL
xlOLPSclCFq/tLY5Y+vUY1EbBUhpV0M4tz+HKE+JJNkeAX72k03cVsdBOeZRlzy3ErVqgQdgPYqD
WPI2HWbUf6KXQYDkNPIQ+6NcK/+SpYO1IOOOETpr1/4Z6qJZQ/t97I587ptgwF5nDOqmkLwaVCRu
lNaSWrMrIYXYqz5FwmOXFOeyfEZ27CexO8nOsevg01RcMZKXHhKWVgh20nh5PNhTBomWybfFMJ/L
VQi1S2eP3RafjpwNbGbPJCeGkK+tYqz6im8x37BK9lzrsRDhMqXjLBzA1XHzE3h4DOnQeaVhwgtf
cG8nDXRju0scYHhnW8AZf8D95uLF7/o5hYIh/8wucY956fDOFOK66sfm94fHHJKlEw2o65jPusRJ
v7VHx3ANW5isBrOJqGHlayZ0V7OjbnvidJDn7QGKG6ig4AZzU0KywrOWsrB+f38Zl8LrZx0jTPfd
MKhBnU9at6ZyBh2ZsXP3iciw9V1VBv4XbxKebipE8rwAaD/yV81MrRWf/MBIm5sc4aPAfn1J5cHX
QRFwWeg9WL6jrlBTjYX8/J4PVwRGSRr7OSIey5jTWefDoS2vuothAYLabkI5xu3MDxZT1D9d5kOX
qmlUk3xAbk+ULLCT3M/aojLdsJPeIptCBB41XcZesQhONkUPTxQf2FqtTXfdUhkWPpPHveNExWf2
Py02/Rt2A3MYHlf/95j0CTcll7+SHo48f5E7uZMDBTehCJGwwLwd/OBy03VCfQaKFwcb7gpFwjFE
lsM8CmQavW5dkXN68ljU2CMA91Z4pCBF5XkAAutpbke5TVvkK2YrLTpL8R3WPYK7GdSZTNF9Tfcv
B00KYJ9HdXEjG+CuYet0RmBQyVZDywoaH1RO/be79yY2XLbBPGglARVmUpJQd+nLljSwksvkxQYD
avWpn34bqCgkw80pn656QiADHD/XkIz7srlqucMQzbx2VRbef7XAI1Eza28noKaUtMBVz8blKSA8
zDYhce98xHxNjDsJj0zKeACVHcmrwUOp5nEDpztLUmzSbWqIvG6tjnROB6kQJyn2/ds1q+kmKszG
1atW+toF6kWDm/w2F8sQ16R2dB0W9eS8Xr8l6G7MxD2sUE5i5yTubS0UQfKGfAtkCpPz5Iphwgnb
IJHqw0BfXU8kZHnk+qGYPlLexEC9ZNEnxWelNCFIDlhmaRD3ZdyxPv1pqgQ+E/z34sH3arZWKs7i
K/9xzMvv+3YEKmcIh5KzIFO3oFdxfYdtFCL07ykJQo+c8xRwfSJ8WcVlZrY3xyZ68VJMkb0yCziF
ZPfM7Wr+OdFDnZ3hZR910u608lKhYs11fCkTbUr8UZnrwoWaGcSZlEMTI8zLTLlm1QEHCwQYUbca
hyYHlgMfWYYdrMfOihYAG05c+N693rHuPRW73WpCUtjgRLd5sU1kOZca/CM+wk2sMFSLl8ikUeZ3
8iXRTMn015QPFgH1jyNEgDdHRXcW1aOft1n7CviJQWJJHO73ib7ZMAWM6z6rBvN1UWgZs8qdHcVs
PCAV6f8tqZiqjeRzYzZtwjCbVpdWrYrqChGdBb5Z7gbgVsR6+9937GsN2y+70p3Y5UArcTsZeL29
GNDYzPt/EaLmffIXfrMMwqCeHWCOreI1Gtgxmjmf57ppA3KrxhNelWd3T4L14vgA2gxxNwFMHjqs
wiAqzieQFD/UVllh/XctAY7n6LHlwTKL+WzUXcRKqaBN0ySwWlaEix6BwnAugp2AMV1v5qSC8ttS
U6yZaacnoH3CyNhnqZE3R+d/B2kPouPYaaeIzFm1g7oEjUNmIkGsKhVoRYct+oheHvW7b8uXl1AS
fiEhWuPaLzSF/cKAJIhjS7vSmVkfq71hDtbOUAG5hFXbjv5Z2PZyfEeWqrK6+HLqc+IFyz8yObqg
ExIx4BwAnObTmg8kjhHvFTgILhz2NNyei8MC/kl3iAkQs2QbWMLq4RTzNq2ePm6ZCD3n/dIqSzRo
IHfrX87PTJxlR1I+dMdV1bqUICx891wcRbpDbzNrzCjn1WangqwKes2wtQi4cKZU3qucFbKjWDz6
tO54fJ6GgAMzd5Dns4Lu6r77c1zacd+FOn/fv7lNqcPWqHXRK+OuFJe+KzrGZwySTVrTYe4BlSnz
Ar+bnHdSeRm7xSQ9b/3YVDxkjSpI3mSdVi9/u9rs7UhDm1qaQh4rzIhv0zzJwbRpDuD50s8hXNf9
QTBAVc06Rn2BU9TfeF9ndAEN34+1tTjae/LuySSwH2ADojuXNhaldhGhd9lV13YZxeO1nTp09Icl
gqBGk9rMnGwt9KVbTSMXS5+QHR7V56kV5pQ0qS40Uuaw8dWDqkZVGDZ/cg/08eQg+xf720PONtm1
6VcJBt+vBWFslQA4osC0Cq4mRJiSnDvq/Q5F7KbrNdUMVdZvuL+nBV6SH4tcPCTAbcVAUeQQnF57
oRJzZ9Re70Zv1wGQx5nNgeDmIMGhaUeUephrVjcncbOgDhIZpzZhNJQtkpuTAS/V+GB4fejNp0Nn
e8Fb9BbBvFMNQUT/zM+HE+nM9nEvIqwCz18JMkqGeCLt5SNzr96x5jVuUs6mj3THGXVcHkaxvJpP
mTwHZhwdSShvJWIc8tzieZUmFEK9KqsLmczIqT1mNov0EnGvM3O4RRizsDOM122iCdH01E4QxJyt
uzQVZxDptSQebz9+Z/Q7VLZR69fbsoGty+6ZNpE1rKRA8pJalM7M5ruouVgK7q8F3dAYVbk+6OHB
HF8UEKOLYQcVyOMbM+XoMugaiPwWjPFLC3cYNqr8EATnVvYiEu8ev3wvfA7+cG6e2GuOZYKFtKir
h//vi0TAxhl0O5kz4bVaLKcKchyZj9lslrn3Jol3bBFqBjS3lWb310XwOkZInFHsZVhcX/G9F/+v
8abAaDfQ5iilAtDN34qCU9iYQIPZubGK9V/eofo6s0yh6FQrO/K2IcDcrP2V+bvGxNvgM3REWqv4
XXu5yOSjnwXstQQF4w1sGzh6LXxjkWzjPs/AwCXwIk0alFVjHlxUc4zDZ4jJsYyuruEQJO0AqoGk
fPtHshkHzL/0bslwiFMUqbhvPIpxocdQrEDD7cKzlO3daIcc2fCvC2m1dAS5DeRmWuaCBxETAhKb
ORve3Jh31nkVY6MqaOG4d8YPHuDhwy54/dhAxS0bVUnpU4wAUfEPVS8YytnYP+xSC+SpRgsfufdL
v0pBqBW2mifCUHhXvzMXKWYAdPikKn0M15W910Zf4d74jOmkjI2QNYkUZ7owUd+xGxLhXk6yWB12
a6hnslAaN3S2J7QiL96I3oNzdRHz7DSNOgGQU2kHZEb3xigLvpXY5SOXTo+93++gxT1K1/tQle+h
0ngxjVR3XttGIXnKV2ZyFTZ3OYLXspjMoxBvA0edA2Lzv2Bqgmln2XoN8GtBi058gvBKjI/CQ0RG
gj4IgBXY+GSb1XtWNM2oiy9swwRaOYFSVTxkseT/eWLjyxK+4IE4fBWQhIvZ04RFLXR6Ym0E6ODt
Q3axwQwZvPHXn7+ppIgC19VQWz5v4MDBriG4kglul65O5LHxO0hJ2O2K2wIMr/FvEV9WX0QL3Job
b4T0yB1gmHoJX5sidUrsWESXZHQ48FY2yljUOQHm8hOmEiRNFCmegpwm50hd44Dx6WV/5NDOgisl
rRDkAfIfiY4+1rVWLDJlHm6l1ENhLD4HC3hSY0dXeCFgPsACoGj93sTNCGOfUxckGkj/cKV449yB
GxgmOzfa1XofuPz/iVeZfEwLLLV9BNV2vw380to6HbG7+35ZhR41Nw0lx7k0/owapWx70R4rjC5q
V42NCk7c3rFpPIWrtEf5BJ7O8u3y/N6LuqHdwAuFvB8WL9QDIGSSMEtzBg/clOAs1HZ7WG+oeLiC
Qd4584J4Ik7+VjpWN2TA43Wv3IWBs28nfT6U1Mels7k/wo010MurVPAXszVyfFyfU/+hDgpJ/mMp
aC9k9IrSbU9KSMflRXXPlWQ1+DKHzrpQWcyJhWOAa28LjoMO6TNRQ0KvMqhahxQ0sKCYqONk6/7A
Bv6lGxZ/GrDNK5+c25e4ny93Adb06Gvf1z4MHwdNdEeJlWGhoG4VZnVU9WkILMaNAkX8t5skadIA
cRYVOU7YbQZtDrmob2kZm1jJBzP8s5z72TfrrjCVcGwU8UmMCs9xXMkqMs8AsYApoxgx5nFIV1Gi
NAQrLEbegB0LPl9WSBs97G52Hgcuo3OV6cfRJh07YtR5vwwc5LzqC3i4r1CUDJcEkJDUbNNNa+X3
1XirPzzXDYwlpUQPoq14SR84eC0zlBaQDcbhl6W67zNT+Z7L2XjDOmDfOi+CqLBMRo4ZjhfIeAWC
B38QNbV8wlxK2ExizMMcJOU91Q5B1by8SJNdv31k1/S+KbR/11HG+dPxzGyFViXbxC55LMjznjBR
xoDH8q3B+kjc8a+RCa82AV1TVsGuKB3hxDo6hErXZsyPaIL7QkwWGBkAHOT3WzKby2JWWOE/GK6w
X2pJo7EhH4ej1FddWOR1fnRlxFitU5oAub6hTxH3gdqqgioeeNwuDwjXbhPJBQ1RR3eew9EQUjbo
AH3gl02kwL23ihQ9mvZcba2ycRbSsOcEvyxervseFLU/cxpP3e+53ypD5/7Gujeh336A1uWDgrjo
jBURicLiVf2Q56kDD0CtCWOFOcnzxZ4AA1fy2+eSPeU7AjWA6KH+Ox9EL3kZNbMIm979gHtEcweY
QSmiMNx8khrvyzorThelEbazRdRvS/WAEHEYS/+Cp7sgV7xsuIqbR21CaiQUaevcxhF9WBZ/hNv/
aufdeeU+qpxou18LOwqgLuvZvX75aoPSGt9/wmjmWhVJ1+JWXWMoX+NcXwf0bCydTG6jRl5AeYm5
y2HqCruPa0rUTQy5powkQthFTN1t4uXsuYCr1GX0H97towZ+QFE3HbtgTx2q1U4ZW2KbrUUSGUSw
6GDcT2sj5ai4Xt0yKDcWuN0aZLmKkUpYM/9DYZC+UDdVKNfExma4UBa/e4UxsM8Zd8+dvVpJDePw
z0EGpuomN+ZQxJHjuyqRuJmV0xuVUZE/tUhSchwfXa501p1vqwP4fqLRwqMUWFIZ0qXyM1rfToZG
TWJ+1xRjdBe8U9H3NHuzkRTqlPSphXKQpjX+keUfaaQIg8u4cJGa66JX3ZUBQl9X9rugObf2YQca
i+s3PIUhmJ7dFfUS4JmwGQheO50SvAwrgaDbTnTRJDWps3MtFuzqTIoHfezEtJHZeXeWtarq6Xp4
b02yTTmhlc6kH6bh8HSzTP44KndCddnqjq7lurqPYi6Ks2kGyNQCedz2o2lUNr8ls31RGXvL1fzb
9Lu2+mQ9ogelC3jzDIlazgbpRCb33Qp+V3J1brIBla22zBSMqvBQnpfogKpj2iq6Do+yM7j9hKvA
H0bHPrCXeXnvcIy7IjSZ9B2XsNvgWXCOPWJY7C3pZmNqRXW82zE6ZdZ2os48+vE/wVBwkYTWW2bz
2idT98nBu+5qRRcg4AaAWZ1Wief3PfAwFyj2eFuspiB/NjU8pBK/yemC5d+wPv8ulq01dWhJ+7Dg
Q3S8xzYW7IvOUgWY1NMppHHaBupZdXrI5uP5xCe91fdzeyjxbksbq/DRmDDBfqhol9391O7el0P7
pKMkDNbJLvTWx3UDgzv6OtyD8qG+WwChGJWnM18zEWwk9l1HHYg+DkptSoUOUI+1mlXX3LqvHRiw
VjddsWPGUC1975fO68FGa+pbxg/34V39U99MOYQQpFfMEy+tRyLQT0dwDdjRk0znNXL9E/tsMKww
+ZD8zB/0rm27l5YgBqw+VJ64LPwHjCZeaDnCj9LHKPxlA8pdt/38oIeDPyf4RcYWFWznSazAwGQn
ikqkIgp9UNkSlMvx7Br66h9uTMN10QPiX9ne0bxcT26Q88XtfNK7/iQNHewvN3ymtNvjllX55vJH
X+uc5pkmloq8x/hwd3AD8/+rNfaggaD3aXO2yEcrFZXUU3+NcelqDlTN6t9Bjm6olwjFGf3llRWS
hIpsAyaWS/oNfovXzUzILRKLj8BcZ8QAc8Zn2T9N987buCmMc8qWGA4Kg56m/iA8FLfNeCQC/kWp
QQ9cQ8GTsfOFHRSZR/9iwWLrs+I3LQMTjk5CLENoKiv825iaYoPBmpXcukD58JGZCUJKMTm7b/hg
+Ssy073rh8Bgd0R3yGysSIQnkCfzOSSBsFE+rZcL4d0PkITi9QdF+yAOeguoQ9FbYistqsJDgXIY
LBumaLHUKrFcCKtXl71FUWGr5W4Z7+omsCTtJ/Rgn4vyE++2Al2cYIJrhFtdbYB5MC5niqw79vfO
14sywALmqeMSkOtkTNakU3q9Rsak6Gn1/AWMfDtYoX+L3K19yI/4aStKgpV5Y0hKrYI7CYQVT1uT
yFt338lJQYsXE4e74TyGxx0fHGcuQ9CBu1IwXbjYbei4QU+gkNcXAKFT4V1kNh/3tjAVqpfTTA9L
vkN421gAv8dGswQXsbBmEpuWMFHrUy+yQAN4RM8r99dRYyg83fV6bCpeNngImxZo+cXBKIK9B2U2
I6IdOyl7Cs8+o4tCiVKXZzQox2S5wsbJD2gOufOnTlWs59tytWyp6+DSXewzW13w8HowK3HMyiT2
YFycH3P2DHbwYPj+x4lE2pCRTjVXfmY49jUkIrG5zTIhxd6j9dVYIM6XJlAVN7fBQ8XJBc4PdNzn
fPgaBSE50e6WQtvw8nVYIaSEGOEcQOCJ5ELuNvre2rk3LXjq0xwZc4R69wNXEI69jbykabJNf67g
Ebf9nYSiJ6zmFTsQdIaua7io3oqVxNx4avN/FF1YDqNfQdD7O9OqlUdOyOhflhDEhoMeZujzWBUw
LWY00cQ1zClCYNAgfss4+oo0iTdK0yAy/ysnS1psVnOwYwV8unlZTCoiDmPZA4u/39GVtMbYcq6P
y+gTxSxNkzkX3IKVvehbhtSx03uNWXXF2eatMkuPADXr59yNy4fJLD1y9OCgEFYuGfyoQtRxF3mg
3Zgo4IpANf2W5qP9Au93B7Ex5mVdhYq2wTqMFN66hpjb9zTCoLSyd9vyPILlJeRZRIxh5Fdn2H0y
zktmOpLHTBqlwYeATBsB1wvGIQVUCKpU1wL/eQSL4Jgmqf39mCuAKZGNRRoyDFId5FUNm4Iv9gBv
iiSXh8x5MWEnnwb1dT9FN1EDxE1l7H73T88nubKZmP+7X2KassaGfMKECrkUjEEb6biKF74EEPzO
MwFKhlLP3tSeTTguZP2shzn8buJ0TQh8KasQaA5sw9v+cXmIGvu7DCDCjKGTCPU+m/u1zkUTNrhy
kMmR7Fvlc8fB2+vGyWY+iCWJ55g+7wnSkB/A35DApLweIZLbqSJXqYIGj0nI9wZwboUsOoXR2cPM
FaUg4h7IY34ngnKgTrUc2lqb8L7nGsW7uFLbiVV/qIcKQDJ2wCs5dmXIRcEU8TsQ6sAMa4kxb8HM
Y208JSmOg2Lq3kyDx6zvxSkTTdrHPxHBd8YBzdMChcOJFH3UqZ2qXLXKbYkUa6LTj5Qi1aDA65Ri
M/uG4FELTN392+JnFLLBNBYEr9CvxMLGZ0UA+eGVtYOKZHBiGOIoYdioebRoI41q9r0Umsl1czfP
alY1Vlnv0gB6IRH8SVDmPN09O8UMELrFLjMNRT+uT3JnvmLm5n+ikEysp9k9yskUPG1Nvh7E1MAg
OvRAsybruqq7b6a2q57YGEBqqZhPXDXeN7J5xsFTYHMT45AKcgwvNAPF6wjhabiPjfVxyjR7TftB
iaG35VteqlDiDTOwzEbw1ICkDf/BNOKYJcA746+lve8N9SKiyOekpLOtdpOmXuXjW3PtDSCiTkZv
puqS88XdEOKxXmIuGHxY59PjOG+mXSFJqFS/IJj0Lw9qa3ZZLOQkhXXethM702myI27kSuWej4Q0
9itKy/3UWkwaabK83ENYTSKRZttKk/O4U14peYKn6gxzZ3KOrL9WrGB6JMYIYYLSQbM2v1l783PM
4k9ofMzEWqmOnwFh4zeKqTm+5DYMCtMTYnTEteYvmEdIyDx+Fk+x/aDLFYNky+xsB7mZ1GahbSZd
uSqyLjbuT8OMInlq47AbAIJ8tpqCp0lOS88/nvGqPMrQUiskowuA+pfQ0SfEyX/Qfl57aIJFXZAI
zqfeEpVLGQqWHiMrg7slTITcRQD4mO3EyTdk0pJRkF9aLRUsJwRdtSM43QAyP41wk6HLWiBr28yj
Uty8KdfNP6XYXZDkjupMlQTXiS1paLmxCqF5oe4E7BaBRiyEGier35SxxmX1a5Thv2XayjPHZ1px
ZzbIHf/NggbvnQi60I3vz7H6pffpkg+4ipkvq3AubwudfYt+x8EgwAsbOH/zAMH9itF8m2oe578b
yi94wLYw8YnxlCjyKB/ofwr7EnzkBV5qDHL7T5r6k9hp9QO5me3YOZJbSP2Qda0s1UFEHa/DEv84
SJQzPAlFhn72PdNo8wozXpW7fWi3nI6Y2U58r+s3e4zReiKgEhBFZwErzgkMTDrGUORp3H7vW18E
75f+wtzH7ZKhr8VBdYeHDsR3R0lZCVCyQfKAeobz+Nfny/ghJtdJ5CZH3QL3QjzeohdLOU9d1ypE
i2jy/+mX22aEmrUNU+GTuBaMSJUWus9jroVGymxKxmGwCvkqIvkusGY3AvW//mYUn2lgdMxTeHSz
xETz/ZU9ecb91x5ieR6w5NtrBSndYenl9N7yNXJSKMPNHu33PpTheZFhenTaAmYgYuHIO6JzdAdo
xwQaLkd4N1jMa0zSrn77HFp9zfP/EH7fEMQi3pNcQmdJcib3DghJq8DD3TdYFvOeiaugj3qjITlL
heZKlzF8wefOgKPbUJUdoPdnqGcShAHcWke7AE5ChvgvcrFCN4QTd+6I7cnhel9JtlEpEpLaHR6Y
PUfMaBQsxuXW+7e0yvPWWinQsJKZCpJ0Yt6/OLVIKKWRWyDDfHkwibivch4LOgNCHLdSMwP4v5FX
Vukbv8Raj1zy2DOddVty0RS7hQlUn/WKLjpMAuPo69g4IBRk+YPvo5rm/D775YpeI/kTuOCyzzMa
7y0cvFkqUG77Qi79QTQ1kXp8yFGSR/g815bmy7ws2jOPTIcbBVKkf0BhXlj13w4Yc2Wuo/TN/6Ho
ut6izMWnmQ//ZECZ+NFotuFkbz6KxPguPQ0+RjS8wNW4XCKW7RzZ9BL853yOQzwbssD1YLi06Nxz
BUgeeE7JI3391yj5BscJPt3Fm1SRJaZnUPq+K13wWkD7H6CeWiP7hjVXKeEHylDRmtRrQSn2PuUF
Swgb6eiMI4jaOOJfr3k47GU3vRfk0fL8OJEltxYwK8+SBgNcj1d25HVUuOSDk/cSFrCXu2/VBAqh
vwMmsknlCycwO/KxCJQjctUiJlE+hXOxbkMBOvV8wSafIrvvYx/98cp91a6uQ5vw/ynpWNrHa5dP
rlXntWdDgnwBoAunG79sVq/geO62XPpZhOPlmUliM9bQIOh9oZhU8pNLD1yl492TJ7gMS8gRq8nT
BW+Bw3armeORcJgsj+zAJCY8kdU0jCtJQhyNMCDmNdVzW83sCKx8xGtpXJTkof5g3udTzcvJqlzM
7Q3+8tFCS2at81WRVojf4KUlg2xnsZE7VIEQ3k9w2JNkRRn5Hx9uV2q/7RV6DLadbSbTaV04tGDT
6yisgMgtb3ecp8jIAgCisOtk8ZcyNe6lCGRlU4ZavcDcvzvMM4ZganDsuDr2zH+nrzeS1s+nt2ZA
x9I9q7zB/b19kfkJOPLg2qxstiGFJPoMrNefr4ISyB5U6Qm0pRtxBQ3TRQbzLbSlkUPJBmhsd4Ub
K8kabXWg8JV46x3pC2uU8ZfGjF1CSy16R49L/pKgqimGulFO/lBEiX7k8CdgOCCp+fnocz9CbYXg
3Bue4ueQkEAbVxbiHW3e1x5LHNIflqfqzokInH+b39TYOAYM8DxgO43jJ1758cxiJEkCifGftGlq
g+LIh80Z+eQDw64cqrWFRVKMxIt2cMbEgC//ChE0GmifzbHI3czs9szpihf7EhBVdezcIoEBok+d
+uT+WUMJEcyxZvVnac3xIQp/FKQGtvPyCY0rkq3AWCSW3uHk46xriUiC0re6WxL217jfDLjN5R71
fFp9dous75Dju+/BiM8nDrQIBAVkL97vEnH5LhmL+Xt9grIZ7wfVxUZ96ynh3cGl3HSmH2XRCymw
1VuE+33WRLZ+sT/weIDyumFNF+UKtVjIdebBDpGQp4L2//fh7IlLsp6NGgstH+68NIy3FOaJyQza
sgYTrG9E9wdlTCwmt9H4SJMzW1vmzV/Nsv5Rnxxb2idXI9lXQcqglvFHP9SviHfbhag8gRWm/ee8
jkVjTqAESW61UoTl6gjH5/1s6wXhEj5qCnUKDw8TwVqtWyeJ2TGdc5bmj70M6vzv9ZSGyzucpG6d
cPuf7ZnHy8lj4m0ec1pf5e0j/0shPWpy1OhEIAVzd8OSO4N92Uo70VDIpg+DHmV7IyLjFEFd80f6
Dnls5p98dhRNnDdlJ3RpEHQubExaDcTZF2ntVtmpazI9B38lphDaVy79Lsxda8nwio7YXZAKnqVe
iFK3qiZ+ZRDEp2qJ1zHNtX7vaJxpMvEl67Vfh461crdn4kUISmueDf+iW/AanFRVCmsshAq7n2NH
ptNBeLCVLXGPkUD3YrZWv8Pgw2Rj4S4mM2MCEYXFSZMGgAaj6S755RkiRKM7t30LdPFNDoY5dZnT
2A/IeA2OJmMi/WMgDsJYhPJA4/V1Ol8iZ7DfyR6ae7MJNsTxPOVLKkKeatVZLLaguAVDZFSNKwop
TeAe7T/UeDlVoHhDHsC34z/3uU8PmWc9W6ibyoKSyspcjXd9VxYZ3oC7lNqssEp+rSWnBQ37gYsV
OHz8Mq76CdSJ8KON8TD9+UOzdTDoX6PMV3+4eZZNKOAPMQogBvDSqtKGTAgTY+rQoCKIUnaLkDqi
I/7pl8mqLdjc8L0KF4i5F5UaFjH+lHwkZ7QCu2RysvPg4AnqZFOMUg5or0Acu5Uslq/df9ZNmzoW
Iox823WwSZvcozovUyKoxYccAe0ss3TfrkE/HlidmC+JWtrRFinYRck2ksM9b1TmJPyUQz9TcReI
uxVCwP5AAa7oMG3/aA6gVLvcWoH/mZncMY+IWQiozw4plFp7k0M7ros5WnRkljryuJ1R4dQfi8Tg
zVZ810/aeOc+TMdxCVtoULj8SRUxFLu1sSlnm/c91U3VWszOU69ECwRntZbLUFU2ZHPjkD6hEvSy
zyLBY08NKHsjutwxvJ6BSOl+tF+xk9X5zGpItsEaxFMr/5VuQggyefU9VyppshYFAf6MO8P5GEyX
4hil0fyOvBwH5oPxu3J1UwXrxA6iYRC8sir14y0DYLfL742e6A2aH+2aT20Qrf7/Dw3GuH/0RGIc
MRQiOOqlB8oXWU86iSL/aUMrCw0ZR5M3ivFFToy9zNyvbw1dxqNXegu/5qN2D8UfuWoxR7yEVUPn
8G8QJX1iTuHaxF7VpGEDky6QYF3+OYoi2rr1UzrWFRovIlXdRTPU0IFXR0DGUuXNUSgQl9QWXdYN
LmTYcqJe0BE8ZqpD7X6UPWkfzoqHXV2jOmlIBRsz4EMNuld3ys66dZ1g8wUYPhDRG+o6FFAQztnp
TWLgAyYuP3Q3jEJ4MuaKf+1+JPZtRN30akKNDSX3I8jHdp5F7R6qB2Hx4v6UKI6Kwuzm3H52vg9t
5NwzDfSQ9j9+bQvJkLrpIcv8IpaJnRxqaCM+s75fvh1dcdQxBQA375sj2KQqWZqQJZhejZemRnAC
DGEY/iXR0a2OOCiiqr1sYtZe566Oj+r54AYTsbnyrzVWnT1Aq4HIQ3fqqK5XkwdHS9/IFbISdqRI
Siw2ITQhvbCyposzGhJtW03hdOIb8mDU053Gd0y3IutzpeJcJRX2P2iK3Oh1AAwnFhZfMLUCz7aS
9Ik6Sv1LaEwT9TGmK4WH86YnnTnI4rTEJNTm7vYwZwwzcxFxOy2bYeDntEOchOAJnKJGgAAn35aP
La/hAL+BBdG4BUx4bQmPny0tjHcYnN/FheYuB3Pk01tqROhnYXC37vkfJF4rOVNCct67In/CFFDN
SqYlCcJCLBT06XnDwo8V9ua33Q8UZpUtFmUoDUYPMvpflssKEJZJnGUD2ftNIL0+tqNncCBMVLJn
+SvOSCCeP67Po3u4ErppeXQrEl9MXML6UeRHJB/KgYAXumQUqUuDdT1vNvNg3lUzfebTV5cfX4kW
zZGXhrYgU8NU86lKDEalmQgtASEisqsU67xGklY2wpp7MR9RnqUZAf0hO0jkmg+OcnHXeJHcvBJF
cD7OZ8PqDxl3lGMCgMN6rOCobP3l5mLr+XmfLMclgfYPAuVYniViH/17ZuqjSJvk7LAA1FF+LR6O
WZhJHkpOM9aVDmOjd02I/J0WHspf8OFrJwQzx0H3bwr8Ii0VL0RrguWl+l70Py3q3Nu8rXtRgcdu
VKtMyjwn0lh03YXsam4P9DIisaaC9psT45KUP7OefHCcQMrdpTWxnEmkSH6bi/WwJSa/r5ml3Z3P
9ClirntwOjMzwCNxrwgELA+DEx5s5OBR4087hqLjuRjkrwHQ3tc/Ob95/vxVCwT/MDkm5vASO8ev
HiEjt/JSpmPu5poMz/dX7EiyBwRpc3IXgPyrOb9qS3ph55rLog3IMrvL8T4A5tnvmd41f9XC9Wi/
ge0F3OUD9Bm5dHmAHYNe/OLpH/hrFAM/ZY0oHZF6oGo6//xliafTJWFl359JCjXclyoy7B/sGTaC
Cj8+51b9tqANKJaGVsAxQrCR/lsA6VnpBu3Yfm9dE2pqwVxPTtaeP+3KM74JmUEG7/jxu6CVA/h7
Evt+m+l7WWVSN7Y9UR0jjJS8YHCvw+pdyAphxOsL5MmZo2qF73G0ub9Jm9o0duFl1JzKX+cba15k
yaBqmrxLgz7rrvITH8auth3bQp5y+N9XtFZ1070DFdeOvssXR8emg3qGEnibDORMdq43KTFdbeEE
Z9XgtrNwgqo5EnW9YSpcGYPhIEJch1btJx7XdbwdvX+9SH9xBaf8VFoLoSSG0mKypq4nyAd8jN0L
PYel7ws49agnZEGNSo4rMXGjgaB8t1rYn5WCF6nq1fVtfiU4J2c03AQDDeTkLcrNA/az+svwUr4e
3KeIhIs1apUrMIu/UhLRz1/P/og0CaBzoehnYuAsTjXbK53vOIuohaPIzjRu2KpTn3kayr3DnY+h
X1APptPg/AEq4kSRxsvFE70MbusQYv4SGNpG89wvdWrGmOLTZa/B6L82vpT7BAUkarcw+JTfKpI1
WJYTKHWY5G+JCxTmGv1QrUaFrrjo7G7kNfolH5H01qDYNA+GLjqSE4qBJg5FeZs/NuQFnMwhccWw
FLoi5yOzWzDdHMMINxkif1GLD/k8CfswL1g+aZZh+I2kGrJspahj6SNoLl5gDBVK00ZNPNyu7xXM
cEkxUUwgoqTLQP6MjItj8gZGLctzrnTdTicnEYIcNEJpyJRRjBveJpKbHbPVVWHmM67ZVKyZCLnL
C6hxe8GRkTKKMudhXNrgDoMfUSBOYj6sPEKbMyodWdud35Pd2pjojIgXblXA2+w92lXoh9DZ4sSc
r7xcAYxiruSxysk2kanYdOXnS+D2fZw/xO/p6lLQ1VE1ecA5Eoceubzed4ideR2wf5rTX4aRrPhd
z1MFAPPuC3M04EIUL1872OPhx+4/jC+8JX5hC7xnLge9LH5p3q9I9AXdFRfQBVmpP1wXiBt2gojZ
6eToYpbm6igGE2rKangyQcTUSMIr/nPE1k3mUTBK4jxPnU0oAriZ17Tg92PX4Q+Tu68RMxSJb+Gk
0ugdjqDqUci2vzhFreeP8t8yFonTuAXqTYxfoC8afs5O3wYrdpqtf2xRsUbhQJkE2rNeFEqxgTzu
VF/nFvflF4bdeNeiwe6uuRn19Y11FT/Cku7GJ7cjnQceXZeL/9LZ7R9PfJGumqcu5J4Dv7Qrf7/A
eC2VGUvoZ/tocBTCbRsnumpW4PMXV3fTXnx6JusciA1o2E7gaDd825Ja5z+/cNIX9k1U/QAkCfFr
Sa5L102ZxTv+UDW1kflT1b3yMJJs0wn+FgFtwidT7v8HOjeJw594DTk9npbajOstupldvNfAEHnQ
nEeB0s0O62EQ+skMXKMAMneO0Yn5JbWiD+XV7xb58lcTQ2epoQVCY/ZVtsM/8sYVjrytbrKK4x5j
zuMhOP3l/RW1pNtq33xp7H4WoqJl3oYMzwIOualUO2gfh3thldvz9l0dOdo5x5iQxD5eHFLXLTaN
jT2WoAV2sk+u5ofUa7QBI92OhL2gxUdB8FRrVDl5BU8WsiPq3affYrFSj6sMMefA73naZuDsWu4J
9FkPraLF5PK6UPSpveQGAjdFrHbgTxk9yi750ST524x5/wrMo/ki1b5c/w0yjb0F0NblUIJhQxiD
ZF/7rlwB8+zpGysoWWzOFc52lqMSr61HegbyFZnM+pUHT6ZHpR57cEiGi9sVt4SJAsGK6JMM56nt
4S3ICHqE5GnQdT2kFk8Vw6V1CwGd2aVb1vLtRPRR/0ZT2uqe0Rbc1i/0E6rY8iC10NO/I5uhASKQ
izK81M5VwKwSQ29g/QV6xwo2om+4m165j1AcTZWNTFijyytm52GPGujno4DCs4/t5T44lU8yVZDD
ifrv52Iio6OIkICFiUpuzvNmKHqmMIEqy1kB/YTUYJXvPOghNVes+OWr3BmJon9V3CN6wN0DtPkQ
YXonpr9muWhD3jkrEI9guYBlJg/2AbZYG72nFF9Qr58mUlvjS3BnK8GSs9xWboW9veKDI+qrexZu
7fsoGBhqGe1XkRTZvy8H6JSOSJfMq0MSG5+y3bJO6encW3+/vezsxkdBQsIhoO8nB5L5iAoZbSQ6
us54RxJZkfVHmvENc1pr1YzgPjcYjvEtv+ofaK1pzVvKN6nufSWJR/pE0jdKlL++ZA21TvBRhqn6
PHFUDNetzHcd9Jvm/xLxld2Dy9wJLTyX/s4e9vP+sw19UX330WMhoXn7qTPnFtSNhCZgTd8xGffh
u3sRjTgTVQXFFtKEk5XlSMhMIloSu6l+xEZroKmXvv+3eAyJA6lfHSp8rcrgSNbUJwaoJLmf5ERJ
+MRXkwbwm6125omuWhOfuKPn0cnEJw0BGcE8YC0+tQoR8dnk5axQeQiB2pmXIVvqn3Cs6Q7JYUJp
XEZ5QLUHv+WjOi47c8SFY93ktPvL6FDpB/eVG/WciX6xQ3W0GUAeknD9IumI4d8DFtTB71VAfCb/
W3t1CnGhKCFEPZ+gxrcazSRSky0CYAhgB3a3jwFIbOAYMvR6n70RwBlXmN4ezwE6pcy8UNjiSSTD
htmZtmk8C12036nFM6RQJGStonigXdV6ghEiaz4ztP0yQsv3E4Hw9VBnBHZQPpABgrBjbNXpJeei
9/aUmawGYybkA/KqrgRWDLPKsfqf3Ahf2mAJhk6nog+N0Zj2pqHUGAWnxSQc4FAG49KufMvieuHI
hg7V0ZXW8xJosGiiSjhdzs9W/wNvALjuxESFj197IELIMl7AHZKi+lPhLSXwIN9Pu9q7LzkXSMlZ
MJ7WJmIRPAUBrtXLBCwTlO0De442Nfe5gWi3D8Ri1MENV1SFXtduzVLTJrNfroqrY+uy4yhh7O5f
bN8w2zdF5tX1x8tRFi1g9/3FkYfQvwly7jtpeJuelt8y7f5+v/fS4e+YO23CrXsZjRhJ0FxSBZ5f
Stbd1LWzu6spbnUCR26iOFsaxhEorfLJNux6qQ3k65T56XsmMa8GtRObaY3VV/QMR59gNrL43D3N
0W7Uyh75VhNnh6PsAs7BSkd+uEwivhclHznaOniXF8G9tPAcMY5k3ojV4313bDNjTI+5iynWWR7A
2mWqsMVPOBqooWf0vmfTjKruXVMKNPO5BmRK5pS5dnVCneISgx3hBFJI8Urc/PJk3LcSbi0KlKuL
kASrh5e41So+/yWBW3ILzbxVKB4cGHboewLyqnZn3pa3c4bwSd8cMy+sNpBcInpurfuH5y9uNrGu
4XPcEtq5wqZusB/ce0QjygGFTeA9EY+On1ySixbCqES6F+0qmkQXHfyRrC8FAayfpG8CMXyHIIWO
w1d0vRcjk8GjwvgRc4s3Cq3weSt8BdsJOMrdEB3TmJzAYR2abo+vd4ihFVjL+hgLn3V/8fDoR2QH
yoR4lgYSUG/Klefu8nfEwpwCXHVHwUr9aTiS/vJjn5nRvmj53QSbl7kewjUI69X/QNMTweLhTrUo
LkfvTb+NzUg5B4+WtAFn4vCtIJFF3qWvlVyxvG0hIsbpVS6hA3hCyua+ku3UHh6+uZcufO7vm1RO
0XqTydO0mkvYTo3qWKko8UB8czo3TNZ1x2x7TsHhOdviUkHxD/hnQOVjyWIxQSBP90bnNXF0s232
AYnagVpZWs002eTbYir59gd++Vz4nQl/A+VbQoM9zCImM1tRUFOwc6l4UXcQ6mnNZxTIk8sEZkSg
qFcXPRCXQ3halmP6YKspQ0wEkCtk5Fg4lRDLHD4ngqTk51vLGQIkCzkUJIn9skA4cbEFcEmWps55
RW0evwrHcF8fIlNO1v415p/3CfM7JdrPyplcw1YW0Z9b7D4i8tERBESHycgMTaCPGi6c6LDDxBNv
v/If9SyxHAegaQEwiUBYD20JQHTpm9ZHJsY8v9sXjCEYIy5OnuWBFWoOvnV1PBdKTsdspb1xpB23
G87n9ung11NKTwkIHTucm0gIcCWzCAhgfb4TadxFxAPsqUmSYKSt7G3CVp5ag7SeHtTEg6ZTSiLE
zfyOktioBXYGdpJSiaWS6AA7IfMQuqJOQJTk0WGeQGe4wAZBjI8n58D1Ma+Wm7RPRZcTkCDsI+Qu
IJkenamqm+p5mbVVM2zIIRSRGhsboiIw9zIDrSp1NZQMVji1AlrjIP3kOLnwd2NagnEd50rdbJeT
L/c5DHSNJd0I+397+qGJJcZWuDJ6ynVBCm7mXxyDVQ82uDG1RbpXCyneJFVMC1SjoWc/u0f3uq7c
Gq6qeoUEOhr+FOisanb5mSJM74/+0WhHz++RDOaKdSvpjUI+Hj/Rl0v732rJMU2PI/L3H4cpcTsk
oVdGJkLBXOZEbikhqXEUFB2n81sTTa+D/tfiKhwQ2uPLjuGL23ojgSKuOIP+R0azyDhq/3wcu2Tc
6eA5G9LIK9pzojuMlSmEhIL2+UDp2IHYjb37IsXZq9fb0rjfeAFsOT4oXbxKuXT3utHrFPG690eI
XY0ND1XrPgWYWYZSCl1vp3QFFYXeBzS6F8BYCSTaSXwCjlVnbow4gFXgTZ2LjqFibg+CA9ETCeKu
sKogLe+fsylD+2AaVAr5SOFW5QwElMllo1V7kue4AFyaKOngJNdRLCFMOMkf/wiCWO16XC8lKaVI
wRX+sH4erTHXsjt6YVeV+1dzzeYsx3YQy+r1o/6rD6uotu7iMon3Wzmdb3NR6LmubKapDGtBThZ2
21YGc/l8h1toCG22WfCuietLYZDQakFYolkohWv4XTwteBDK+KeKzn3OurGb1p4aeYuzNJkOQdD1
ohG+XQt6d1YlfQl/4ckN4FNGQARyDeA/RsVx4ioUtof9HbEZgrQR+VnTv0CjaebEuoxUe6lbbZLe
3QuNfPujxs6kkY+pXzIUEowV8GOxMD49KoOOweUT094hWB+EdFaBkg9Fa2oqmweevH4szFJzh8a+
IuGIQUVzsUwUSFfPeD8AZm1sQrUZZcjvGvA5Dz7db3QN5GxjwEfTwm6CMoK5IcKvfXUjgzrZnRgW
UyWGDYj7J0UhgBgnqS6GXUOEQ/mqdkuxMH90jBHJKxRNIyXGewwWYLpVRp2WB7RxceVAmC95nll2
8CmICJwNnRkuhleOHglymmn2nbIfAPZ0Pg2IcESP3FjPDLiovRbMc5NILQ8e7ng8WxOUczsW7Ank
Idi2fa/bq0BFhVoHxOOXmBv8GiuWofv3jIZ23otNbyAL3Mgp6eDc2C95O0vGyhRn8UKPmM3Bwl+2
qzQoGid1AfLzsviu3ToeeUPq9miWnIi7DPylzzqQPkxCORpt8LLK9z7PT7SRy+1p5yw1HGopITRf
EvjRzrtj5AsamcmV5n947wS8Vz4bj9gJy05T7rwoaUs87U9AVot4XuVjPNkmxcNE0sKjqbtw6+8L
7g7g98Y62vE28O8VSPvapfXSaSld/mGZJKkDQeotm+KhVjYD2WilEKLTOtAL8s+AGEdhph+WpCJy
Ps53TpvH6toJEDyYf3le8UQSULL6W1HMDeTuGHeUSeAS3a/iepSwhauXxiHjT+96Heth71JjZquz
xnclAcxS4AxxvAUBIvtwkRJqSi/kiFZU5m/wzYGX3LTizVdwYSi64FvV7FO+BZWVG66719/93K2p
TLb4cocqD5qTTfU09fsxSrqYBWATWuekLjWD7cwtiO3PbgZ0gg5d8uwXPh37/arlfyKagZMjGoFs
EmI5gbIMtpTPD/Qf5uKLIT2Qxr8Q1S6Qf67ZgM4LIv0pxEI5ZU1N3zLKSZHPC8h8V3SqprFUDSDW
20Lk41XXo9Ignj0t8nmV1R2wxsem6nnjrGxyR0W2evIt8WLJDDQaJiLd2tVphLwzTr01TSUCeOJs
XIX3LQ7otbkpxW/gYmlbf0W9gguDYTkKvEIUKqoWyFiO+2w/DbbX1qst0gRsuHG7SbX8NKdx0wfZ
Hi1JXjCZCQaOOzjou9SpYpXRNA3tjl5ijwlijuXJD8cAxsGdzmwl8qxJdK2QBpuN+zcTBpRSvlR5
T3FalOOSl9ThdELEAF857iYs8dereyklhkVKnRdreO9TntRTvs9fbeReytVBbdJq0jDQ3PTFrBnB
9BYnM3mhtn/GopWh767SFV08opH0kI/wboeWJ26bC+ZUqs1UBxJ4OUeaJLci5+r7zpEHrxpXWPmc
xjGD51u+vjZ4np0yGIJRq6YwWApMtoByELB7A/aAFced1ilZpWNMgkYZ/Le8Tf0Qc4z0LULkiQkL
T2pqkMWG44QkFSAzxvY0mJ86BX2ERMaJyKEQbGSakAYpvV51BAmUVHpgIchAXdv8NEDx3DOCzA0Q
ZbpqEU722yFTQiecS5DSMBCSYYBDDk28sj12WG3tUPkeuK7XQjeH47DUG5YytOeiBY1RN24bP5Px
5xTjPLaup6E88ii+Cz7Ii0RyE4yFJ9UTfk6H7gUIn4JSCGm/lLmyr7GqlX2VXjcrXpRUR9BHl7yP
4HZkyOrfT78Pe01gViGmuRqc24ebifHFTIksjWyzt1ILLW4k0KxVD0QI2TgiJxm3n/jZkg/5jIpM
x6hjjLDU66FNz8maC69+kiY3z7pR/JYd4KeD1f+Hf6mCXb9PsWQchgB6EWkyeQ52dEZfqv4olKYy
eF3usFu+ueOy6132EX8MDJ3qA46eWFnaTkng/7d3QHU9wZ/T3uSFB5i3ZpEWLm/2+VsZa67+1aks
EXVExn//j5JwgcVgg59h/s5I84xDYOs3XTShWDzdj87WeEcnZIZ5jJ3+o0IuMsWrjEOLT007gHes
Zspyls38vTuIaxbL2P+TjdlS5JbwLvmYcSMRewhomIfvbgKitA8fLxbHsCwzAAjJFOkrEk+3293A
Tbg13SlWxm1fut4Syz4SVPSU+nXhvuyCae+RBW23YUe6IA2W7KwnJTW4aTqrtKfvyi85yq3Bhju6
V3Nh/5sH+oqX62rTrhYS/k6SZiuuxSOcHKp5PFseBM8pYesKrZNs/NKCivs47+Ns0dJqHYciqlWv
SRf+p4fooZ0S3RKIgc8Zcfv3PJPEB5L8GxVF9Iwinym1S8UHuY+WCnsdRNTF9Z5A7+DpV1AJBe99
7ayr3a06bUsEwuDVSkKp3FNOtDVY3QwGqArAN7fnVL6HzDB9xi48bLCd8ap4jrx8U2C7BXNZYl6w
q8JRjiuIRqWymItfqwzoFSpromzavHSApk5MLg23JXYgwv5NIz7pDn4S0kt9Zq4iw6PMcTR+aTct
EslEZt588i9meMqq19htGFuctMsYCVkSxkGnLsO8Ks0e2qlwiyA+J1NWAuf3dc9Zgf8DDx50sn5j
Q1oXQ1uqXsj+6HcDGB77c9P7QBDewd8+bQoJgeoiMIJ36rA5ISX312eFlK6ix5MTytBJ+ySp5dt0
evq4pNLAatJ9ZepHGPEhlj1Ubp6A4kmLYZMuXBuoP+Dqj4wL0D0mZh0aQaEgddk2qMk86cP03fbe
NRAVRIx/+KhCQ2No1qRE77UktXfxjVax3vJ8Vl3tPKXu3We6SsLhSDWMGeCogO0qy91YzSENzMMv
1Bk7OFNcHTNf7nKo6slLpnodWm8d6jQl048u8OHeXHChlySkT2/8YEKt7x4hId4OkJmnWgju/PXH
gMBde7ypNeiek7gLE4/BZ/BW70dj2xVqelsHVtgimKiagb2cKFUj5PnJFgwLREhJk/7/ulckex8H
S1eDHxq+DSPCfxUozc9WXLduV/KBSoHf6dt+f5Pk0jycWSNNYxmceIXeQzqQQ1C1u/FuWQhLmKRa
WatDvmpdY8RtlIrxAVv4BKp/pkPnTVmGeyitv38/QQTh8Mm9t2CbyLdtCZ+E9Q+gDs+j8+ZMYuFr
prfM5c7TxWjUN0CrE2ko2aEHyCIAuxYLy8g2lXGOTrz2Yu9EAlhrEIavIx/KzL0DyXrMr7SKHAYH
OlH6vUB1Y5r1O6i4pfHNVWy6byz7fK2xAJnGcAf+QCugZJoZxjmh8Y/wR4xlchs/yfkQQLUTN5qV
yRuqIuyWgTE3XlkseBGgww0T6/hYs9Yb7tvIq1Q8WwQZtKvZrAM8pVlSNeHE7IoJE+Xr0RTU7joi
yCldF6F5VQaDU1c81NLcKX6LlSR1DoTxQMvlMEW2RHbzQ0ZmyPejiR1qqTUNRcZ62GrfkVhwNocH
xoLW8HOE4YxNYoe8Oz9yq1ciZIK6kCTI2NHWm8/u6dXA42nHmvHgBbesNtFU5rFQw+okghbu9dmH
wYqzPVHat6FP6rlSa4ejPZFdx1KuTpW60ma4ysFaWEuZbKTIaj0tmRhqhnMpP3IBmaQ/b/1R/PiC
LQ7KLowSvCCNUTOMRbjPWFLgXVhCjh3FDkLV5a0WqVxzHlt4kE165XpdIaJvSC1uBmpAXGuenbWI
6kWg8CcgPiACTni6mId396zKHhYj6K/Z+1QlC+Gaur9l5jP5ohDLV3v9i21Fp2af/qWzr3zjg5T9
CJR65uw1RbllZHD51lxH9eFH3xfYm6jV0hQyBxwCORLZetxOvCI9gz2H3+lnvUESHu3GV3787IzD
hgsZY2QPhvisx3b19NspV12P2CcvHQcsqIcz7TJKx2peuzehBdPCT0AJ+Fvxmr9GRgepVfav5Ils
a0mDVnHKDLtBKEwekFvgU+fRzsYgn8plT96TU6SifLNxLQHqtWmyONogferXsjY6R88GtsgWtx3b
/YB/W7l10L/WG0Z1lpJstbXnSJ28KMfs/yCGRHrbPqli7pYnN8J0tW+H+Jj4ES6OrFJaw387rVuv
Ehb2+abknF1ZybHoVxdqDqTfyb9DVl7/YIR9cV7jJAvX/SWu3w+aGHzVvVw1isQVoMVRoQzuaOyB
E095I8uMjWT78c5zzWEO0KRcH/2yT7NFXm1V4n0Tk7UFfh2NeVHz5iZoddqtHefbIPAYP++YdsuF
os+Axbenk+FDOMK8LuChka+qz+UkH5o1iS+Skysh2sNEAiWHGwCOIM21SNB/EDNpPAULuPUZaEe9
CXjuKWxaVzZjAjkU5B1rul7v7FlOVp0f76ZEboCmsMz7cR27+Q9ZDWYaLZHKRu1lDj2rIjNA88rc
yNhYAsBqvMznYq/fKXFU+McWdV0PY6y2ut2ZAtnb/p5TnHdHhVwGl3+hop3WR9VbOuW0Uk+FOEMJ
QHClXukTBTEeL69SSy3+pGQKc4myk311/VcpFy0YDRzCizZ0UfHU41reXZxsE5b/Pr0UOKhxWaQL
OOOW3xsyinNbukgVArvbfuuQk3xRmwnb1bgvEOKssbMV5NL/N6sdcvbvoq5HTW/WhRos7IA209Fz
Hs2C1HmlmJA1cDDclwk9Z9wxYB+o7d7hNkMKFRFTRVgkpoCKjRsZALhCjMlvjay5P3H7wCHZMK3/
GrhpdA/A1sDa9eqUl3+n+2SJA1v7jhlpAsFyq6p7C1Df9hP7PLTG6CsZ+cevYCut70yvHwKUpFKP
rbFHzPmYg9C6M+4dtieai58loLsuvBtuTQSV2/+1sA1+/edY9WL7mLp6kGYDR2HVfPt/FfMmF4sj
GwoakQ8QgMiiDXfiIdStKuUXUaUAGfUH28jDtBN16DX/7TFEgYd5pYAQdu42eCqZTyaHWQk9VZgi
C8//UTTaQjYncCVrkIZJTlXABnqJsh5n5DJ8dRGZL1OtS+ARh5N9oalqiDLDirISU05xaPURVNOS
jGFm7cjw3lQhHLleQHEIIZNFv5IksWTTiOvFYXZxiZL2c7gOq5Orv3mGa7CukFQNOgdoHADaI3Ul
+hiNnJDj2nxB1URlsJU0lIvpy67ls+5s/wAbEqM4APnOKAhy3l+aDI6vrAQRLVnbZRHQrw4x0XYX
/ZscEm1Y42En4mbAGiIIRvBQ3Auzt6lZzBSHw4Yl5PQ3/fEg8l0nPHSiW4o118cUbSxhRDWwCsDr
oQIFnhR/vsez5VtB5sydau83RqQau6YqRGJcrHOASoFmnl5UdxRPDQCE9fmcf7JsWZHja+4pcSXT
gGSRiQUquZWNm90/PC9K578EIBgEgCVy+oOfFboBDM/Pdgp3hBVBkXOoJYC4paP+R5M8exROi+19
HGlIV2fRzoHJyhcH6naf3XwCK7ecbZVznnqllsVanFNFuUJJWbaGvfhsMADwu9kSqMSaVMu3zzdZ
5g/4CXOW5sAYS2WdtJ5OGw5LoCNPShT+tQoKDcf6TWy19N/yMo8VXz6kJwfLaFwKXA5pvJWdFoK8
rYNvc1GRhZ7gR3tPbYwdn/U53xymJvLmx5EHYmXdM3U2+lKbMPEaQ35RSPN039jEnbZ7wMLu4FMW
IuqwA70Zu6zEX5RFqPYqPZgITVpg3aoEzZnRIxJeQHdiKt2YuuiWmJv/VkpzZpnKknFuIo5+IB0/
RnogyZMmBJqa3BMqjCiJR9Yj7I5/p9qw+jAcMrT3TcOa6dh3Ohb2O9Z7G6mTxQyr30bESnUXI2Ks
OMqLi/oIkv+9lX5Jp3tWW76QZLnvtjlsB723VC+0eU+NTj/vbQLnMhtRWyfGk9blKAfiexgeD9w4
4PP9Fiuj10sfjjN1umSfKKRusQ4efT7U7Chu30SNnFwM1Pdo/SK92Dtz5hKTj7uURh8KRm3menMF
SFEosXnwg3zioQ7NbYgUTpyYZDhCE99f1RBTl+O3E9YrzeJMUzIMVg7LrpbYLt4Wmyg95Xgml51f
CT+cWPuWgrDb4YWk780yiXYmS/5er8DOZgilQHfo/X5WVxHghfOXcfHNHq00448vIlE8FJ8RuXuo
ucgUcjKvVHEUS/wu2akhd1Yz/UDAYRlvrIDEv2B/6oKDKPZdEQuUwACeDTbaCtwHKqkn9kxfaaoQ
Wqj3tVt1EOV2YIrCPd0hLAAGr4/KkkVI9zncS6eUQ051z9JtngSW+qolKvcSWhL9D6HgM0VKxqzU
1GzzeHF5cSuW+4wMXBVHWIyGgUgQUoXP0g7yfM8K9FWO/X9wYD7F+BDTLPoKU+Jh3l9Zg8zlGM0U
gXUd1WeHNQobuYTV7eiAc3ikTLzBRxAn+rplY9rUfNfAn1JkZXjj+5+lCPBzKaRw1XP469qlesAH
qyJAFgd8GYj7b6GO1lIQTyha2iX+0q9GBRAWEAZ7l4Rhhb7LT+wDKMbL8fyMFasPbkm/Juz2Ph7p
EVbN9A/INWKPRj9EsfHhZk4668CobF4lETjG8gHEkz0u+/uGOher52QkD2Bvt8RYJIw5mU2er0r1
BkJ468YyECEFTDNLhntpOhAiNjplsLl+vx7MFiO5xsMNBrn8yvrfnUKRs5TbimEjT4l5VSH3tVQi
h2lqHw2Pj41yLzShu6pg2GNz18jWkyVj2+6+7L4iMOuJ0YfOcDn990du3fgM1upbdwT0mBwYU+tT
YOKsyXsodvmVT59ptR1M25tblqevvICmaXC5ClYnEnNP7lCrHChugmSE7PnGHZVPQmlwrPsnWCl8
aOSLeSkMuQHXvDJGII2zCZ0zsjJTYstsdfreZoXbI7WFGWCKnPYsV54XX16szSBr8q0gHDkdXpDJ
PnePIxhnPLreV3OQxlwAay++R7x+++XYYTRWxLGf8GlL67jdcZaPORswVcAxf3cTIi4LHPDwxGEV
RXWQQ5E1dSBoJbmrf2Ph2mTvTOOY53YrzOqsZuBhHG/ItAt2f4MR9slHV9kZXVDpdLhnXLWpWitl
KrMqj1IXMEm479i10UBNZFg5aOE96e3XKS7adeXIqI4Wez5QeP5btkV4UdTERNyUF/Mw144r82os
uGtRvEfSFNnmXgy9LZx+EkC7rBoth/jNtrWEWpWyxEBcVy2Xu3oQz+khaq3iOpVWJo/ZXxhlB2UE
EGCpMPfqAStfP8rND/iBb++kfZqa/rNvrVDb4vLJilo+CmV2LSy5Sbg4hskM/8wAttih/sYt+iJ6
rWyIKzwD41UZ+QtaTtbVWNhZldtKTIy0gep0HX/dh6brGkz7E4etmKOzn4cRD4DE71kuJkaPxcMJ
e+mCHRy26Jje86d+Ewr4fl8bIbblEbjBcAdgp8S5bM9pxq2w4Zhngc4zVlpd2qiwRuQwmnl+Z8K9
7liGimTlMFrO8SCm4e3pZQsL79qUCiu6MH+1DTLB+534XGqGEPym5aFBWEz/jtbhH/oJf72/cogL
0PG5s/rJcplpMExxxAf8VVoXMNJJ+aSqMxNORCJ3gPBGYWnUTObL6JtEmGk4tV0WdagFhMntDi+B
F6aHdlE8G/AtM6mgHblrLssTQTf9StVdFM1pZbeeEKwMCOZQfID76C4XOGWVZeDWYWsHqKBDNPOG
3czJCouU0VOIsIbEQIZNxLE5MrkTXcY5VN2drbh/m99b3pLbyqGpx1LaSErozOuiMDT0Dh7ZyIjc
WTg7D29AZWhNyZK//UyanUCGA280auvS1VzEM7Pgm81vg4QxYqhcx84MOWz6qdyUs/pRTTFT8weJ
U+lV0r0OFfM8yNVT075G1F5qYjwHfGjyTuT86CfmbxrtGw3QlWDmSMF1F8czCThoXWqya6J6181i
cGMi41OQc6GM/D2Aap0VbmXqsNmnmxPPJ6WPXd7U5xwcObUdnfM8BUt7HBQ++JAdImGZuFAfFfe5
ijdO5HJYWWmP6z/ZX+IgAdUImSmf60pYeptspOorW2xt5zfX3RbuWef8KXFcBJhgHu93MPkFtMcQ
Abk5FTnX9Q3uLjS9/3WN9ydUHAD1ynN4LawVt2EUht3GsxZ2JoS1lb/K1EgsLPptj7BU3yjEMnzx
CsjLtS/EcF99JNvyQR8qn8lXeSfYCnvdXK/AtTS1zkNmIFDRa86jOSh1bvamUjqWn/Z3ch1GVLIT
O+dBrvZwmS7CjnpTiRJV1dwImfEiE97Gcjhs/oBhU77W+48oTH52VYvV5CnfoGSbmu3xr8yV6PgP
ClvABbiI0d2N05CXBCr86Yau9GQaCPsXWaVTgyQEpr5xa6svVg4rQcApReicn6q10uJ6CJYgdfFB
0MWEhUECNDhQaDmyOBGJVjbQUaa4F4SF4sX1XyTn+U13CAenUdSSIjk0Z1nQnTz0BllvrxLULFbm
Um+9lxfKXhbjXVyfl2morkTU2VuhMzm6C+JEiH4X/gYEXmkhcqY1fUSF/zFaEm2iENsJ73p2w1eV
jBcs9afKXFwE6TpUftEiQr4KVI+Hp65DX+l7w7QpwsbGfmBlFLEefvz3sJjmDIZWLFHqEvkXV/od
/nRRvZNigyw6w7tJA7EB6xZUiG6ZkwIcGC7FaNU2TKBOFvyLTixub+j2ccFQFEQP1TI8BGax5bG9
aDg29xnj7MCZ08H0BqrrY9HK7Z8+cKEthkiYmkb11TYcacqWHMf+z8C+BbjJifTpktsOyn4k+RU7
L9IHefMUzLg7VTv7hu3zkfwrIeOg4lDmSiTYiihuW94xNNLjSaBhIPQjkjHPDSK7jrSR2wHEl/M+
oUgHkxktYSo89cr+r0GXuLDL0ee4CwnDd9jvNiyMB4z6/bG+qZCS+esQNeLXmq9JRRzIRlUWTqgZ
4fqO3M3+jW5G6zDFVhLsSKAFPsmJGVIwq++Lt+SDXDPvdeaWFhggRF/t95XPdNlSQZkJPTgm9hWM
N268PRwv6CB3uauZ6IxauWwIhB2PM10WK26a4NBCXP8DR2B1VynqTbhVydJjLp8pyueieupqc13M
XfwEF33CmM40idBeuztyuEJ1WciZPD7N+FCJn+jycyDsWt0KEOyM7rx/TxsLHCbGXd7tEM1my27Y
KURlVxaM+Gdp/SbUc6lk0xXm1sIicWXMa71rlvjdOQi927nCCJj5vQzCGP+pD4xT/56kLx4bnyf9
+OACmdiNjbWN9wl+lZFXw5olG/t2S0N4Rhipnu/iGoW6bHfj7gbkoN4hKMPf6bDNNG8LVcyirPCg
6Hu2nbNMe4gXDt16Gy7RFSDOgDROo5iWGaHD9YbYNi0pF5059dCOka7RuEP1D8rhWohgfWavddi0
EVUvTrsSFfL23Cjp0paepvJaOCyGSZixzU3Gjvl6Yeeh6QQBwIoz/5qMVoQ4YhzwcLwA5F5zGHbQ
T4ic2HaHem6Ak2HQCv6krtTalrZsxlykaz+vYFB0bngOXSKDxCQfFADucKty8CSCXPen4txJqsI0
/HLkHazcrDk2XTPcA7zqx5f8WBkp2XL7u4gPwyWyMOr/eEqvnlDbs5+qq6zJuzTx73Sh7q3t/lVg
wZjXJHmE+gTVJBBSkb9mpQ7+K+o82V3CxhofzefSzOYYj//6WyxOyk3e+b08gih6XL7Bep+oxTjk
zgDVFvAdowwIbCPk11kJaJgz+f438JALUwNnf5Hhk+Cm/IzA1wicHfE3sdruw7WvXmesIOv9fg0j
Bc500jXs/n0KSU1Ou120OoefmeBwzAwu9jv1D5QOLfcRfTZPbuXdKWKgYpct+wBAFotQVZKO5w/J
f47mEZ8eXm4i7nWtuFLh1YjlMfwPOHh3ixiL9g/X0boyqli4inpTIBXfojXUSI0fJSnTBMhFoDfv
P1DtBJET2rOunr9pxdiegQublVuneP4AvGinoA2oDi32j0kAjXxAF+SrvZ363/010ueqebJ8nl47
MouKE6Up98ACy8maa5+KT+FaoNAViAANeedOu2vaGOhvLRu6boN6yCyENYEZ8u4/KicIv+KwHCM9
WiugkATwXNV2XouhPDvB9G54yVFwaywINrqjWUOoEpjbJ/64fY4oUcTebquXlsA+O8Z5dTlgT5aY
7i80+/TDLLotsv5cRdbLJz68MtkG24eZXp/onGqiaSz0cw0G7qNB4ubLcid2LuNz80hKtJEQfZiO
BmuyUHFf5hraHDnKO9b+GeO5C27uNBMTy6ug0rEeKgpZcMAl0/M8t0pvuW9U88kg/2YC1LhkxVO+
mLdjIe3zp1SE3QdwAVeVynNfvCIqF09yKYFiLCpoN5XE3H76VZ+7kpARZgDPnC71bxgPUYZtIyis
CQJiOxOWboJ70VhDXrVBSsVHzoD6YI3uRcbdRqrXRAttqvf2QBeKtG1I3G/ENx5nUW2HiVHM8tPR
oSQzbNqkL+dpjzxvwHeQbLaHFsBF9OF6JX8vZLvccP+L85rQCYe7ezD2eEA3/4L/1tkfDnX9fIV7
6p49glT1eR9HFLKPLtuKQywerFyrLvDcO9vEbFaYdG/bPH5OFpOtHwGRmdys9KEtthZdi8n5oZHn
k83qorHhq+FaX92wAQGlsI/EFlxF2MwtNaGUYZvzK8BCXABc3nB7hLfgXGxWUOc+mM44kGQ6wrHF
gQ9QcKmopGKTeq/AUKwrT04a4QJncbemM2LXsJQb/R2RZLpae9Ik/Jw+SLJqrtgreM8lO90R6Wte
G9Zis+qxavcRCMvj4/LXFsQXUlBFS/fsLf5RcGc0hbKPddAo8jqQU+VIP2QMtkwRpM5iEkYihbFa
fkCqI51eTLPE5VnCLQMQhOHJ4RhS/8E9MuR3B29UmJE2XaK5jjVU/4fqvqD+DsBQQYkMVT0d5ir5
cGcaTNO82XCP32AHwm6ULc/nPCW4NofK7w+HnwXGMnf46IMJzt/RUrsU03X8TKqrgcGc09AvwDy3
DSx0QEwVZ8aKXdl1huvxPs8DS0V7hUKPiuidw3kw9qe3T+jWGCpp1UQPchB31Qif287i9UVaoX4n
TqtjGIRE2TL9DHGuyBXF2jQm/r5CvB+qvqp+51vC9LVY+E3t6GU4KgCchrChKztnHzVf8d+CHgkB
dHKF+ilNL9KhME5qtOfRXMSP1ChDpujEfLPx1PbSdsKVxZAW2299hr8uv0zSvGewvzrHSAeNDbZS
+vXK/04bItsYQ7Y2w5NhFuy72U5ZZqKO9yY5dpAKWZZx1RDG4xFazvTJA7bfqLrDuGHKA17FMWAo
9346rAyfduxI3kMDqblCbhUELeQm8nx26ErY916NkoDkgGpfJi2HpFVEYN/F/4vU3pwxyDD3zV/z
jFUdFlfDVbmTHT6QdPD5MhdMqvI3zzTZxvGgiIowd5DxGg777Mii7dROf8oQ1u/0vQLdqx5vQesP
AGczWRizhxwsEhhfUrwtq68pQ6fn7PPKqTZrtj9UyPH2YMvSHu/kobA4ttvhdvv2woIFoz5Vkynv
o4EzxqclyywPlIUlX6GdTVrqOUMuVbynNpbyWcO6iBy9KtL/uBXimGMenepb5LabBIcqE/2jUJFH
17nZUNmehYLvyZeF/SmH/omi6XtqpQkx56l0xNYCym8Vv/F8zU9BkJF+KAfJU912cFikZZDRGziE
1QiAHERNLQxzgAlT2pvACbWOGUteLPhOmJDv+szGBnVzykermrWhLA8Tl3hOE29kaPQzuv3FIlB/
ybRH3cuQCz7aQx25CDQ4BTaigXrDAIGRxXCTzkzlbM3cmG1o7RDkPvSPcy6DoQa3G3gEl8HLV0f1
RiaP8VMfTpT211hqPUJRyYSf+q+8boMnK439olXshi3W4Fkhd4iIUELDsGxwd09KMFdSlKmR4gIt
/xbsUtuPeDqXZHwEmlxwzI5EdwWxLB7tIMzcwsTJy/gAHLmnFh/ptODkEgDEtfPdv0EJFwegU4im
/sTkLsGS953WJePq6Ol2nCeP40QYXXKEazC0KNDDQsd83LXm1zGVrkqSO5j77KqhnxdONP/uykf1
+gDz8fxCFCo1sbSySDPBL8IuJSlhTrJH/UJuciSPkEBizFg22r3qWTQ3tA4pbylhFlpfthT/MO+m
AVACRYn+08HSgmg3l9ycUdZfbleEp6UkvCQPto0ywlIrpVke1WNaGUzocIaCWOVeVYHQ2sJyKA2A
zPfPUTiARtcDECRkqyJdphO8ZoXpZYuxM6EXfe+gvTdCF21C9L5MNqMxXgoXLbwQ3icQYpBbMu2X
s7KJ1dFoEXDWUK/qRS5AUvviZaJR4f7A5rPnjV9UIJQZZob1p6VCtzQpSGhWVIn5kmYEUFDc/Lmv
ndfoAo9DvpmnNyIyZjRWEJ5CQEGcAC9aKJirCFpqzfK/r5N6EH3+uCkdUwEIa//tQnyPQB4Mgfi3
RxST949lErtAkRezukfv4DlNTrEKGTrQEPh24QQRwZxSyo9454tRrxwmFqkFTzmvCfPL6n1oVANm
DdBANfKX+uacybVzJ1gZ9Nwk3IjawDNdQdmx46nqCep3IhE4szgTrY16zkZ13xCvQN/aRGA6DoH4
zJUpWFnRoDAIfWw+W/Vpc2Hrq8lOS0fdK9yo+DOOP05eONCuw+y6lagkDucsd6laIAGBKWkVqy80
kWMOFpTUjzVSGIWLS0+KNjejIwXZGmbCwtxt40e9VLQXQ66BAjbTtaTLxqQnO2hmD9pCBVV3GNvg
rmtw/VpvBrFjLEuJc5dEwjWokrsJFYtsVAKoM5jqz8RQCr9hTQ40lpsG7x3q0pw5+hAd+aAHVTIo
nv6Mv4xVVPpH7gpQy7DOLkBHkx8+gx6jvrSBAPnvKiCwCgD+x/8VPlBfpnuNm/HgbJ1GkUDavY2j
vq7Ul7AsoAKOwbYgpRVEGBZINwA0+flbx4jxRhKYPnaif8Os7kw8+0hefGpl9hc60SY34CcADteJ
xwYPTosRo7VLgk1NC5jVWRKa3O+X4VrYUN6ou7w0pmWEplVv8+MHYZzu3H5K7oInrLh6lQm509nR
P7HpSWKkzjvOHrPW6tIr/TfUigdLZny4hSQo4WIvWRntaMJ3yvLeEiOXPy9N2VWA13ffWM0v/6PT
HDbu4S4IbLT/8gZmNGKsfbRXJ1Fq5TNQI2v4Bqea8+MJZaPRzRnw8guVEV8W0sWFrCMJm/puXBrO
dV4W1ZMoET+1KgYyPZGaiubMfYQ+7x5Xml5DDnlF0FhzY+a7oa68zTOajDN8HYq1uTFk5CcrMi/Q
/Xh8jcur1DOZo50wR0JzbJdVaxNqYen9jQ3jueXNKk6rsX8cLfhSFn6TUEtSami+kWsYWufWWF43
KM5VIAqprzLaalpm+0jL+3EX5xfijQPlnBmnWLV80d61KhuDhSl4/iHQmqbq5tXpAN1HCAmGCG9P
OoCtNr4thCt3iaYCoa0EZ5i2294WNubnXLNi9RKRtbCVSHmtrQ18Y7g0/dipWdDunCwe05SD3XNx
hIaQ/BVP1q3U62WwDgKdeRdtzoja7zg5bx21ybiDibkU7MgnhM+5TmoPhV0E2siGo+gQ4cNio66s
i7FxYmy6nzhVGlMKxafRupfz3aKeoIlNo4/wp4v54530feWZNexCK0rLvBCF0OExARG15DqK0aS8
gv5DgyR+4JVGgPHqALw1cDE81m8EJ5wuf/B59oZ8oTfNyQrHpmgxAvERbXpGSjBqANX1gk5tY8DM
0ZjmZoeC1q18OcgmlvqzSWJ7lQgZu0eMcwPKaOElrZ21zjYgIIYSwrqmWO6+woC7HizaGQLg5PFW
8mySSy2my2iaNHyqF5sMAWgRdS/B+k7edbiGIQO86De+tLO/tmWVsN8DORZqgrwuxyRkMb3ae8B5
pmPjBczvpv8uVkhtpb1IWZIAZDJSc+7HzlgSAktqRCK/hbJfaRm5tn+WG3rIPPn6TZM0ca8r2HXy
WhVA1Jqx5lapZ+OmdP6jM7kh6VSom8oMTq92qk2Mlvg0/0FjCJYgiJ1YKlCqJDshgJmQrOjcQN11
fXxBlhGHsD+UWOwDNubrDUmcGO+4J3B2/WYoQoL1f+cyLAPPSFxfbjsz/K2q6r1tHchXEAfQ5Z6X
VjL2lXYY0FUppw2WFS/4S/SvjcbWydugTkbWvvtmoXuriE0j9uTMoOivst2toHXBf+8PchJM1hCu
3wK2tlsffFrKZO06uxpObS6TAtWwu6tE8lNGnxLJ1uAi6lmVK9FEkBD0I+83+5eK+94CEMTp8Zof
fWmW4LPQufM8G1sozc9PK/Og2HudfVhJLbgQoqWvTqU5jTD+GqzPJ/zG68d27TDTBYjImU0mJbsv
5XoCEbowBOIembSe09l97CCLtrXNxazOB/AsZhdk1/q0z9uV8RT2BqzgndjJHHVgLXwRAVIVpoUh
LpQfXvRIBJ8gtvC/d7jPVa7yXRH8qxEK5yjZMSzQSehTDRVg00zJ7jy44VnAPwCWXCh+CnMlvSQa
ozpZ7fZkpoAiAoiD9rE0X4NPbx85PUeXsvcu9qc0HG+jRjW0JQHuO+F2jK0Mg7GfR724+XoMwOv3
iX48wzYGqqN0aYEd5iYohnZbvh9ToANQb+bHn0VfMz2/eT3X6KOTHka6ROy8Sa6x0QEIZBWqS6i8
wlFaQK5IHv0Ddv5heBVx90+T/KkukNxirWAO76xXhBSKuB5ndM/g6TfMAa5Ss+5la2aIPrNfC1q1
i9DxFPRCnyBgCO7Si+XyeQpfRZjZZNJ8fvg8fj8ewLNh9iMR7n8CruWtxx9w4w0tpw72QyyzTMUf
yRkS6ZUpzyqcg+9MO+wFgp3PgPWP5tuVwL7kyGtFUfk9nKl3vxeBtyfKLl6LmPre+xuV/Z8Z5Og0
MPQlWHTCPiEckcxZ7TiSWuyqaCTYUiM/R7cCoCGyE6MZX2V1LmJNQxIfbs1HzeafXDCkNLI+FQZy
6PwkOz3WlbO0AbjiB0EZJK9iU0KGeNf7dyZ2cjWpaA0Su1BRzl/KhHBSsKjmRO7/uPv0cguBEyDS
M4Sp7gqsKMTsyoSPKj5ATPkuEC27mUMeubeLiRebWTmHEhS76eB4W/8sqTztDJ6Gw23aqvLwwQgY
Fqz8OxSMNQhYQz8uID89QXtfzrb9Ia0MecpvuvEaGPqGMNATkZ73Nnb3HYLHlYfKipwd+iZDNL0I
1Fn+j3hV7SQ/d2WgV4i7z0AE6bd9Vko0Z/NyqFOHnzzs+7HwAeINYwGdtdc5TUCfdz5VghXg6PIA
AKRSLtTIUgy3OPukWQyJL+Mbd5jz2iDqJLiwQH4zww1mFpRkR8TvxQ001Cy9Ai/46jdA3d5nfH0O
R9MQ060P75uzhU+z25OyoXpcmH8s0fFTYJaUYSyhIxT58E1FgBGOLWXtURM6m28RRoo2prRxZwDI
GPYo5R40C60NiJZqdMBmyvLM3qFPNoTLlKtEJz2D0vQEK0IF2hNmD5HvnOvIDNaQQFTb2cvs/OOv
G0ngv4808yF7Pu7NREAgB4AgaXFPx6VzBLxQ4A43z8ur8P5H6OR1QnDBYB4dd2dQpx296xXFGXtP
k/hfgTRDw4D4CQh/GPyM28m4wchIXBS2c5QoIgo431HSt6LZZiplpE2wAko3L+Ek8KDsuv9Y8u9l
0KnlnyfHGZ4HNVbRSpPKCWSxo6mcfNZkulk/5NDVOXa9g3J0Xv58nyOlsRB3H9v3xt2butYSH1VL
DZSElW3u9OUCgc9iO6+XElIGiZJbARTcyfN9eds09I/nSf4tQCEUhye3vvAMK5jJN+EpRcZv0Jw1
M89qauFs/PkkIfCvTYtiV1f8xFfHEHhm+exvhJbLMITQu9bzI4JKi1vs3bqw0yYPymJGHpJY6jqr
4kB874aWOZmdmwdlgDzPxVy0LpV9sIoBeHQeC54eVstJFIIvM4G7tGmhxTqWreDHtT0onO/nRzCs
5YugAnJxLZ7vEXF7ugn1381bWoJoOKY8ohaTevQeTDzkY8u4b1TsP6fENMhlny23ykreEefUpIxZ
vScbQXjWrhz2cFcctjQeyCBXqpOrE/RW0wVG3C/Z+Nmw3MuMP6MljIXxKmmDqhX47JTgo7SSrAcg
kdB7X+NgapqYQOf9HtGM1RUfZb+XJhXt4R/jmCRinwMClyBpG3HavK2o6bjsKCnzI0ONh8LtGL5B
Ic8VahCM6q1VjvZsEkxds/AHmkcuX80ui1qXwkTLxaAr/paydUkYMbrMgI5CFc//fegOOnWj+xmX
Kr2McGX2iAEtnp5RZ5KJ5qrHl6LDE3vMEa87MfnNFusOahI11TiihLPy1qqA2X5DLH+ccIjmQ7O0
MS56HdVbugfmjUABUHJpW80w/wYoo+3zhC0ro5p/lJQwOMXcEKAPc2LqTep7ChCKZXv6Aj+Hcl7T
UJexdBEUpPXgtXdf66467AuosSkwiNJ0xUch6gF6Q6sIsCnx739xJiYjOe1IwWnVneVuigvMRk8L
J4wIl9Shf8vqOaOULYUEN7xX/poYvyHT88c5wuI7XFWLRw5rDGTGa62CiowC6Lsjp/YshOzRgzND
ZKIZW97S4qhDeaqktX1HZRGPNzFJ6Y/a2b382N6AUHA5HDFbGnNv/rQsgTbjtl4YmK+YXzmbev6y
p9PJXBwA0B22kW9IQ4VHrdv//WGf1Vca83pjjmmNoMpahzE7pntUQexo8120VfxIi1nuCKt4+NBV
PCMYRSaY1fYb/kc1rEqyOQ7UqbjyAHws+lYlaxn52YZlxgr277GakhF2uOExTn5dQ9pafV7jm0/0
vptn+KkcCAvSvlIpIAKPEJeiqLuJSe/lFllYdE2H657gzEHCiJhnJxQebOWTqhc5wRF4gs6KPoXb
pHFX4kCHMPGwp77Lg9zaQ9lotVqttJz94+q3Cv2+kUW46Kc6W4VIhCD2YR4aTyeeYrmxYpr6uKnP
iqdU6a4eb+C7sCDpsReSH13vO0hKeF4mytdegJlJUciM3PKhQtejz0Jr4/xcI2/iiM67TjSgc95k
5d50YwrYkDynPfGouu0vR4gceUJVNeMWBBiFrjo9N9t76xNAFYC9bkoDJ84VUyMDLeDwtvloq2/Z
LHuedoTblK/pLvgikArrPAkpD1wOddQLbRZbWOMHXByL5j6t7Xw7W7L5AsiB00CJCAtwC4mYKAET
dRBr9vYbd/72V7BlcWsLZ2c4RB8eSmICJK5xHKxz9FbTPB6icLpdY2ItE3X8ZDxmmJJCutkj5cnt
XLemJSmSGJQaZ8Gxy3e1fkvV9enGr/q9E5CEFZpE+VqwesBvI+irTe/pqSjUnUBSdaSNV8Nrxx5W
plebZcnYSLqnXHR2fJPyKtQAJJ8a9lfmyQ3lYELW5Q21PPubQSrSn4pqA7LkjIY2WGaYeNkRVTwf
z8kB0sYE4Jh5q0J/hCCfdjsCN35/oMKjoG1aQWSzd3dDYM9Q+u64nDvQt2tkXZAj5J/9TAsw5g4e
vIOsXEUeD7d331t1JbJlMYeionJvtXLREnZTgfVQriqrpLxF1C+TcihXy7A6QWSwwvBPwz1SKfRP
rDqWnTZzcPbgcv9GNpOMxt6Kt13o/SjdMWW1V4Xe9jtlqY3jfCYNXtKtGtKcZUl5wbO/cWIVgzeS
FnlTpP8A6uY2loBI5a9P9mLJQNeY/vbzM0uZiysaovDyE1iXlhYFdE5uVDso70OJMZmGky95VDvv
drlVAf26p7Zta7rEzM/zIE990bILgP6HZgI7lMcIvcw/GknCuW9cS8IpEZdcUJjA6Tl18WnIZRjx
OXzoI4bGFj+f2+mvjQUUbzAfdGegyv+KTHI910iofQbzxAOfaHbJ+DnIZEWWgyZD4MBJFx5fMSAI
cI643cGZiFcq9Z5noQNDGuUQG/pBR8/hNPF+u2x2ijJ+/t51t+B6COFxO9/YDvGuV2rsukzlkW+L
LO1pDGNKKDlTgjj/phrJvW5AG/9B5zt/A8xKGW2SulJmFzobJHowXhZjEWf+kLf6QiNBMtSSWtZS
K36uV9cWAq54i21ZATKJqOmNjkkn6lPd4qiVKMPteV34phXSV/Ln3h9BQd1eo1vCu7/waXeOeoHk
g+PcWF8mg88mgv6UZfdxmpQG6jgk3yobzQNyMdFBTLjJHKbWvyQUI2Y46g1j87L2MFALS6pJxUOh
NYHtTKoLu4MHmN1owReew0Asfp282KM3b/rghiyY9uYP7EGnPdQJ4PWnt2S+ZintYt+NVBAvzODO
djlypb2+PDik39qRgU09TVlWu8qJlyKRebmAOmJUwMZVhK/R6LIxqVTCNzn9oeRSg6bUbbBJ5VtI
G8jXnRxCSrS+TI6djD0SXN7oM2p6FkAtOvRqG+a5Zz31tCqe9PPEj92ce7Rz1o34YcngvDmRiRbL
fv8Uqx/nrgHWBCGwdF9/XWbPcmKcz+xtoB/IQRkTW8O8CrDEIGzMatLRCw8WmeN0ZHPQWTQ36f7d
m7urw9+5y7IlZXQhQld9QLzna1PsXWiG+fH+IOD1Q+aldgHMAkfVExAkaRsPmpQWa6HPaeuQmbfg
RU6qec6T0diLXJ8o/C53l+lauDmzEqMEcupAVMEHR3ozqhiIL+BaQhMr5JooGccDD/UQd14rNJeH
l/tbqNdnEPobkDSWY95fUL35fM8uINE61Gl8WHFDizs6XxLpUrWw3eN++qebWKVozv9ur/nih0ag
U4mRdFaB/tnq9D+dQHw10qBLeOibqBgllR7cqoNsT7kw3ISG0ezzFZov7YJfpdBSd5AGgdvlfAfh
mNGCEzMgkLadOctgGoXUUBSfbfJTcsrZrRnFcWIdhy0CDzMX8PJ++NeZI4c4FFOlek/micNfOF9h
bW/3ES+WuQLc6kjmf6g1CtmNVcHwA5NK4ltZxau8rUtch8DtgFoYU/zmPuA8CG2ZhOtSlYvAUxOy
RK7G2QerH99gj5yQrgkQ4Tgk3isuODjVJJ5RUVhoU+oHR7vP1YGLKxVCQgJyOHym1ovCuf7D6ICN
WXbVoH/nZGdJKm5U/emAverJb6bRpJuFFfYagTyOaxVXrbEUK6HMoQficJxmWbZ55ygUTcaQQ22r
0/dDlgMlPifDahaS4Ff4TR72hC94MM95xAPkcz1p3muBHRRNkHBk6CxR7WsIuS0Ffd53ZhfP5ykF
sA+6kLtr9Uspkf/2MdiEDIUaDVZ/GWlAJMZi6L0GMEIsMJin49LM2DJYJKb4tst0fI1JIuK/e/zX
R+VkInAgEcamWbwFLXJSAZilTmccJeCGxT+XlHmpQgwNKJkzXW10zgOK1fvgSxj1Hms0QBgbGOxM
5f5m6MP/+VeNiS3WS2hDXftZgqIjMSZskaNKktfdX+8yosdMhdwks/B3PjtuFrlQHz3cdVpB3777
56b1gGY7hvqwOG5zsFjdaVh51N7QITbgea9RkXGJdM5+ObtXBU3PPb5hWBagFZX1wtEalXZrDSFE
8C+DPnASyZC/SVX6EpJMvtaRjvOfKJi4dvz3iIpIs3383Zow0EQ1PnkNhUJBIIOqpD4Zu3QIUJ6c
Mx2wtbgcb4b8ZW8kuWOeHTouYp95uBqwHDO2mz4KRAnkGIHFN1ryXACSpIpm5S97qTIj1Z7m9Dei
lkW9xV7c0NMzwMgH9fhIinyHe94gD/jBZ5ENQKzBYAluxT5ez8PN8sAgx+lbupj/nTcXXLpILchH
rVW4sBp3TAjq1+SO8HIwDxr/1maF/1CHMszlC+EYjHPvE+uisrxUB94viieEVyrPgaqFnXFBP+SL
NGvbGHmyv6yfZiM2mKYDjz1vIML4YE9BaHTuTSOBfUyDxwxLHJhvoBs8j6zVOiv4M+N5mhXhxfAp
w/DW/1xJILu3XWi38asn7aG6NAO7/vMpEayVlf4RVoqLUMIiZKVxksioKjLmyFJrD+y7e3xKDhJ8
zOda1QoNjLof4R2VexhIVeUNdFB/r/aqNcOt2+pcDVo+Tw87sWoAmdXBy0iJnnSdgo6tjqq2QNpL
1VLrgyvFtJe3nwa7K8p5O3EvBLKTLEscCSrlI1f5aEIYCjRIWUWolO2OGdjiFFwYfco91qxEUh/g
MVHeVDdvToGH4RS/PQNWJ3kB+KvwrzkjDsVhs2F9mTgkjsePEgs9K+xcHUq+qbEu94Sz/mS+DxLl
+Op/zGaYiH4gloctbXpYih9sZJpQgzX1cpBdgtKYEXLQQR1QA347Hrkrt4PD9UKhqm5xwBgrvXgz
zjSyspERjQoDcphVuqTxdomkmTDVPaYOsLr1xkkhZc7NRxtBEKEY3K+rtrXZpPLpAlnazq8lPsP8
NszQqJpQq5raKoDMFFLFltFEahhn2+bu45VbTMr5FP8BgSGtk2gRIeBjfV6hdfwRZBFzqbXR0M/P
GisnJ/zmh5/ElnBDyH29UQeAzPFxPDrbhNjz5Oaos0Se1ypdQ8c0hOCmy+o+/JgDdYzF2AC9JgNa
CSVsPXxc6AuSA6cW0J7k1FSosYOuCcBCHQ1nnW+yv65ITG92pa2ArAefAZ1mmbatIRpssfBpKABL
9ZS3B/dYBVPVOfJT8wW4VZZDgdROTVwzDtJ8ta6xwz/IjgjIeqiQnI6i7s64CN9hvBKCuUCBNuXS
/Nrjet1TzKk5unRJEUir7l/eNbJ8t11LQng+1WLD1IaZvbz7GTh8saYLfhIlYN4c1r5kIYYkcHvY
WaUreR/AEOytRcCF5bQKeN96qTKMFLyB8D0ezOHPaV6koDqQ3SjMhByopIqrW7pG7W3Zl4B5CWpD
3FS0FU/aI6YNwUV910+GVXKQSFLVwTdALFRVZRPDLXmErC5l+Y8ULiywmHwxfys4hY0OCnhgfQLT
7mj0vGpuOKak1+KGAQqWzE/4jnZGbFKuOsPT7t6PhMN3Kr7r5/n3vvyTuHEZGlOaU8vLYIo+Iylf
3GxpPjVwhIrzEm4ITfrD9eieL5WWRWVNMdV0m8Y5GzyF4+tyS+R1bOZw31KKjfEMAURMlu/kLtAy
oVDRTwkXlziIpwgyreHHdoVwV1Lul+V8EsnSo/QP6J04gzvCxLKz0Pqb7qeSKKlShTEo+IN4PGN5
bmbbangWf5l7PgfxquODzOgbwNPSNuK9Tjhjx+C6wMJPLWmAVhVZD7W2WRmg6HG2iAipYOS8VaR4
R36SPWbFIPoAlo5pw5mlw+A831MXGPvjWAvuRmje4Cy3z7L2FeSChwGe0xuq/kmH7CLwIoIzff3g
+kdGf+5VEvM3ZZAmV9azFzHt3WOIdHc2/HJT64dE1EbDHaukDZNt6HAwQq48/S08aFA6VDr7HReO
RZ+V57s93L1beyKrU2uzQAXZKnjrNC3q5JrXDKhyY815Q9l2xoblBAf0NC9fHKyS6HjlywkgGG7v
ib728PFGufWVkXMdTZiscgJA+NaPXWUKqwcY6teT5DGDyYRRicGfrOH9nkBAosntB/WXnHskO4W8
XQCOgolGmsoVxcyfRp/MpXEUi+BmhbfbcxMvR787kLJUEemin3ZqFp/b6DcrvjOA14IER1xovhnp
1sem2NlHS7ltnkVjjsP1DFleuFHw8ZCwcPm8sZ893N+ZIfUGyjAhWfwiowYDEWUW5PH5CTQCay86
G2oE+4K8T4am/Wl+KEaqOPqQtuJP5LC/QHhjBEJ3za7FIQsF1XSwA17aH6oOJVMiY5N+cgY/6PKF
mOxM67Z+HYm39EMVoyFXbxX052NQ9ZZmZyM0A01Cv/8dVAp4bLgq+IIMylpdOeVE2VzWxI3QiVGS
pipPlDHOPeT+o5at7bRxfpyE/d9W+eSFSyq41AdvQ1SK99zA4C3MctDYjh/VPG3T77zsi5emJQRV
IkTuL99OVQr5TjBh68ugDEWTnj7k4qbSczpE6zofi42xZURWW3KQsySPd//8NPK4rSozjEXZV4/w
2uM6nDuJwKBff97KX0kE5Eil57xVQErIpP9igwd1S/O9qaLdprP/6s4vELCX507/4hw07eY09TAP
93qjGQ5GLGRvqAsR6+avc4ZtG3YGsNjtexrofKvDQe3L5bw5dL8jPHw33HOOfL+MwBEJ/k+4bu+D
12gXloCUW9I3usEXqgXNhVTBy8RK5u3Nd2QycteCjSFJs8OBwtEb8x+Bm+GgM0t9DP3yTju5BK63
up3T6XUtPRF0rnwgOG6scTUs6nBddu/pN5Q/QBH2eVzM7tYG7+quO8Y3gDf8hswywvG+dzX/f2od
lGFg62iSDo+820OoXL7d5ZlEP+UAutCLDLxAi4+dzitYB71k4AqWErl8e0P/z6bUKDlnjB1jNJXF
Szio3bh0xSVYCLA4CUsMc00cwc5F++AyVEk6XctnnOeVJaOeBC/SMpl7tL6ZmhLoiq5buUIs2vNk
csRN9qDXlEOtNjvblovgKIdbn3KvRX6BItaob8azVWA7nbi4Uiv0c0qwbmROvHPVtL38E/Zf+91T
HQyoZ3C0w0abWXyDbehTbH0hwgm9xwhKvPxcmWDpaxhzTqz8tzwVPMm9Wxm3KQo19gurI+yU2r1W
xg/NY/oZkHfpwctxVgI+GSKhBXh05QXrM1RzHDt47tcpzByim4WYF1vDM8+3K7bLt4rViYiXbPko
VPGxT6d6l6mHrfrhUHV/QOKNhKrL9y9QZNM/ucRJOPSjO9oGtfmdNnnuyYDsY+mK7ruMQEQiV1Ye
AJtGaMLYXjZlU5s27eq5Ylukwqa1bdhy6qSei89HJ91ma8/+a4xPWfmHKT+MeKD6GFyEeJ2q2Gnw
SZ8etkOfHFWk2j1RS+Q6y2YBxEbPMpchq7twhxUasNF7fyi/rUH/JTp4mY0+7+9Re6FsDriHqfjp
IuyKIk9uWSCrqbFFBi09VPL4jG6rOxGXWx5QFgnfltbij0bNBwr6tlhp36hQTxrio7YkoRe+CkKS
naJbBleYKgltcHEtoIRZsFSoZHHeJt+M10IFZXyAQu+/m8V0sZ9TmYJMDXooqoaTlc4jEJZzQlxm
w+oJOCUJjQxM9b1o3tEjLBuFnNJyu/0wSO1Y4RvG/URbt/IXXtN623ay6dGWID5JykkhzXzRqLP3
2Rm0HUQOpk9N0m/O4FXvLPeYHzDnNO/3xo10ENVhhGJoaduVH/nRc+24skg6Q7um9VLp/z4GJIkS
XUHjEivCedeeN60fFZPv7vsCXFuwWm91gHpSdqnvAUazZUlVd/qu2ESHygVobSz/r9yEa5ay044E
iNBCF7+jZ1+1YCwHMa5xmv1EInO6gShyfC5DTv0qa1i7nuuPfgYXOpl5aW1PpNGG7kPdlURnL0bv
IhdjFNUdghh+6Q8Vz55koU5Vea7+zxT3A1/bqiKKbS5YSJwNMSVzQAC5ylkeEZYVcFyhiaeRy7nt
S2334RdiVhrLcq2LQ0fHEiAYjkBbrdaywPXQkhbSbNMdVhDLmVIV1CwSFvF1kjXpSDFmJrHlw/hS
9SS6UI+lorksTabhAPksly8n9XUMp1m02n/d9Tq+6sHDV3+73ZJp2l4A9FYsovb6pUnGgR9YlM2H
sMU7dNEDhFsep6TO4WEDPvuQuBA5/xY44VtMkE0DKjutdNr1KsECuRc3LBH0fAQZC3L7C7RtrfDY
7xGfymxoIrNKdiGT3wHm3x/L/dGxxrwMsqHUSaY6H1EI/4pxewGCeWOx5qJJ5iOs0lqSICFOToga
ddhEleLI2GbZ2F4m+bCTintXYoHh2JeIzFXzVkc3phvS2iKXUlfP3eO4O7faNiS6d5E74AAnbNQ+
Y8t37bY++sH9qBFbLq6irizNKgyPpYrxTl8M78pKkWKiYdxORDflgPHqfMx+MKqy6aUvBtIUshHI
ltdPy/Ke9OjjphetAqiptFbNyx9XC5Ws/ZSt0MfYsoCHRhkvGt7MSkNsRd10l6Y+NScTTyDC8uX7
9DcVcZMzIKuGTfIzOExjru6yD6uq0qxAOxPZlihoMjuqH8lwEeHnturXyOuXaMADFIsoGfUQmO5n
6skM7pdNpvKeV897tLn1/iPp7yNVrAZ2d9DFZz78/dFBXvFTFfKPmKqZglFxFwOkgjd39ClW95AL
/jjJ9IyWT5lwAX1OvC9k9Vc5djQaJMQ9Kola47Z8Uh0B3M44wb6eN6yP7zQ+sgqNT9IeifYBVxTi
1i7iG3C1N6SXVLQrwHa6TmHBM+VV5/OnqhiX1xUf2iJBcXKlxFOtU2lYaZJdLyvzXn+urC3VqXq/
MVAdayNjfquGbpdCDpt31NhAHIDvBjJPv1mdupAup1yHQxtDQt1CI/i9soNgrqtB1QQddD2xCDI1
jYtws+dRQQT0n2BwioSSevYk+Fg7Rr+bIUj2OJryPuXDfL675nZ5NhiuCtlq7ZjyS7xHeRGrXo7Z
nVRgcp8riOIYSxQaybw+UjdLsbjAbV/IigzLxTvVhjdju2YiJVVc56A6cOattN8Mwv13Uv+DGVLn
g25HOZPZEcDteWtOhmvNfrQZRcLlbLCT30sbiAJdy2h92Wkat/0vCFAfa6n0AOxYsMV9A0Ex3P8z
6DUX4uh89BjRsMssDvjtxFlGgUKO1eA5SoxFOk4UQhVfAQQAlZw9OUqtWNkf78NWh86DTmixtwnj
zz4xbacKcqAP+sV3dNQYfSgjoeaWZ8yPuLFS64rsxNAzIKvr3YkUv0DOFePVL3IHJ1In21DcWZgZ
NCknbK2dhsivE6N8knsGWNTfrsOk6kLUaWoQZMkc486oKrUhyVdYN+rD1vv/XemHA503DcqKEDNt
ugAu/xmxIYovf4v38EYdoYtqqHl3ZEK/ajPs05+a9WqKgZUZvuCslnHZpu17Ou72FHIQR2ASVFhZ
clH95Drqz0LXHKRhpM0HYpPGswY5M2MGsfLGd7hNyWHaFCvtF/4aRLwDe+M5s6ubAXtAVdp9sDvt
o8/S60lH0NQAZ2uIycPJGuK4TW3At7CWyOijzzNttiCKT60Dxq2FkWOVxvwbojEOwK4oo/K26hdX
qc6z/TbnErGfVREWmVBEGjrxEIEGCeHmAFNtT4oMopa/r0BCgPfAQ+wYFFdI9TGf5Y8yLqf2HjGY
K+6zmXTlNQlhdJFhCT6AjSvD0laI3fEBoQq+F4SA/rqV85FdlBIuc+YdMhsd2c/B2REqV2vNLAiw
b536ZU37KZj5RVK1ylVtdyc0Fv+2u0MghEVbUqmalZhvyZdOZam4ru4JpbULJ2mTXCU9STZdnrFI
Szby3hV081Zj+og1aBWmOaaMeKIJEt0mQGzX+GFLvto/qAEThU84hJ1YYNTJS0kx8pgpu9TxMR11
pbl9KOfo2OijwMzxvQwrFmbnzLcaG1gFbkfRGhHI2txaNIBonBtu3Hn1JkcQJKROPmN0QBJBaFnq
tIsG+YcF9HXpqteCeFC5thE+xIO7vn5eEcHMmdcnUxT1RJpmbgQzDGaYorhEsWWoKTjrJUrX8T0A
+7M287pKCcA6H0lZw0lXqQgPQ0ZegSOb+HY4pjfBBSD/R8l7LQqRuqZpE+MrngGvTqwogLuo2hnx
HOS5gKNwXKuLhNxIwUUrV7mh8Tpyxe6InbHgUX1dwhi8xGXditKXqUC09Y3kjH60bsfQubg2ybcn
vh24ld+Zf/S0tyBzdGN0XcLp0nBbk06WwbDpxNHJGlGa68aD+4PBa+ClOsecStzwJq1Me6HCe2Zq
cuuHw8KKhXfOStPouKCgkdPLD/JePbeggY1ZTdOQe7qNrHTSbFWzxIRdpLGoHB9bsvD2bLakqo9G
rh8Z3mVkfslZoHyei9sG0sbAJvcKMcB8FOjdnPwcvFr3rWuQfIPBnEt17nmbrffp/mNpYW4Q124A
1tiOxfVoH2axf1oA131+TSusUISztRiGF3BAU32S6SKK894Mir4Tt8Li5U+6lV0tCESI8fAZurkj
x9/JhTx5RJyb2Gnqbv6GHv/bcdfyC36v56DfTdZ1p4DHd6G0tXRh+glw7DNqjM2WiAkTk066lrzw
jDooHL7PM+ta08xf9/QZ+5l56QoOL0cNiYipSj4rYkEbwYOW4UR5vOWtxE8I1cuF5XccyZW+V3j7
QX7zkpfFJnkAuB/uLYzuug6f9hOQNau7nHRMxfsl5krPND/fByCqhuNrLqYpkKL7otgthPImj+Xc
v8gzRrUlCDhLcgHphDeZKKCXONNARxN9NpOdJhIQaboqlUfdldg6wWl+oLH1YxtyfoHFxoh5p8YX
AgoCuLG3F6b2/HoXa2oTlUUJwOcX0X6MRuyiiqVdoPcH1kQu22OKh2Q5f0buFgao83IoTbKEsIbt
0H6IPe36FQTWIpYAaGAAFowN3hGe042bVIBmZKGbjtsGFX1iysxJ1kFvdakead45AtTvCfezhAYD
jPDVsUdgv8UtUBTnbCTnrDBujpwCDvl0UC1el6J+b0O3O+NotvbEDGpR9W7qcQLPaNCHnNcq102g
BWlT1WbfDGHbBBMf/kgcWrSIsuk7fh/PlpHJeyV+xtr0VIewH2EGgp95UUp/V39g3X+qwvqZCOJl
00LziSI8yb9GUB1HgSgQLu0dPGFczxX0tr5v7TF1iIGXN6WATWz66PROZlah1Oa5Wq8io9CpGAzt
YVsyiwz9+tXrE8f5//14TC1OtaPr+Y5FaUCFeNJ9ufDa9qcDGdD8GlkD6mzJmDCpmB/etd2t/ULo
aIxy3h3VJBNTCs9zoNz0QnNjaMQ/DWYhoA+JWTB1fr/lKY6kOO/RmEn4YABuVdIipDo4L848UgBr
l4RqJgU0O4NUqdc4Y9C8WyqHDDaY3a2oQ2k/Y94vJ/AU0Xc1Zy85xNp7O2YyNUfnUXRGuBlyi+BV
Ej5mHVk07+ZKmqUTKA66A7/sx0PTTbbMYwfemCPy9m+LJEvED6jEiqK7fw6Gfb9w61IGIR0BQHtR
/hFi+9fVqdC546wg4MQzDHUEYNh7rjIv8ZOAKbNBUCJ4b8PKkzs3PYm7svbP2huB1fxV9IIyRddX
jNNnnL2pSQH7/hgBj8BbCMuwG5kvsQGC4bPGSNH7ciDrPL8Stc6P3ptPAWoUeI5M1qfjjg0edYa0
iURo80mDLWnF+BKWSZTICvd1X3tZ9x/+TFaWTEUNxbMZ+556I9af83rDepghKdn32sYiOh8jZ3fA
CpqktldN+Q4tTxNbdHeOJ6gSFCqFJG3wYeNZ5idIbt8mifK57xZSkdirCaKz/BDElio8dK6/2+uO
zqtPj4fSUn+wGF02N33tkb/0FTOgPRsZwCtfQ25nY69OPIQXp52nhrCwx5geXYuv4JtUHtonHNto
mmdsKwaTT3IWOIeEq4Is6rJuo6IYdNIPiR3q71XyVme04K7px0gIvqG7cC1thhQqJ/qfTuMgbbFS
absr3hlpKPoHm85YJ0L0F3/8UXU4SkYDYwyrtZe4GBMsaSCVvyOtcdIZHrmDY8XHjkbO8GMPiKjh
OVt65IrTTokEr4axkB1U64gLjAW7tweeQ1A8JDOYawWeIM5gw/09+3tOxu/+N0/E6n5BTBCOFcba
V6ycuAEjYZEOw303ipT/HM+mFPVxIjxK4LHgNvrGY3o7y/xoZdSfMrTtr77sFyBxaQOt2ppTRAta
halcUPryGotq5CFu8B87DvK3AJ71ksokY7mzuWgkowMh8zH92dCfbNn6ENw9s5GhcSj20HkG4oMj
IDTzlH1rZKft7wvSl65PRku26/yZt5u4u2H6utppKxE/wT8dN1M+haw3kZdaTWQbnvQoXBHUcp6l
J3jaU7eZ6DkUqVg2zfrZ39Fuxld5LXvNr8ac2lNqL3DUHziyRYZrtLwx/sSd3hzq+ELg3ed52CQP
3kmq35PpxRbQm9wDQd35CPMXvsPWDWbYMpeC5Pe/OOjdsW7v/0mc/Ydr5Cf4b0OYTTuj5NIw9DL5
HRDA9fYZEkwzhHLnBTe3gK+3LAzB38EBmrcfAwbockavWjyS0LK4hkOoUGoHu9sbI0VDpz5aCY/h
dGbQzc5MUZBJDrpNwHzal23wywkPquLn5j8AJ7prEUUmTOQcr1mU+uGM1h11PJir9ALL97NqbHf8
q4yNOqOFRYKb4x1BegcaGy+iCep1OmSClilrVoqTEAiH4RR3mpQfUrG56urBdujPhoYL6CYAS57n
VrWKSXAOGIE0wnk2OSthk1De9mxCt8fV3fTBze+oGlEmuikHT5Yvtkky99a4AX1Iz1WrEDqBkq+n
pE4XR5APLEkGWo6payQRtnZFpyK0XF93nhqZSNTgaolohO0u+TKPGLgRxxLtrBkUGIetAtbvIEBq
KBnn3n2Vk3o8KoU356KV2KcbfjwyUVAdH71XntQWBIB8hk+xMxdrkV3/slyWUkX7qXjW3bdM8jZs
ZlyUM0LSwcNbNf8knXO0TwOcu2w7l/NkxanmZHIB/Cb/qu7yTAYQqtg0L7jipN7S10euY7aeWTN2
C484PO2DJsx4sJY4VYE8sX7XdZx71GcgPEVSjiJxvUL13AoEWf4vZK42cgWpzySgzgh7O5gFZl8M
qh5dQLpoRJ7gQagMfKtgwKrh9JX5cKciKyHvnPPa0krImqBgMtEJrA9iDy8lN6xXQBaw8hdKV6F5
+s9230wcfm7s0016KaHkjyU9qJSRvpy2X1YWLuBurBF6UnTSXBj8EjXYjcU4O8OeMf4aW2Doe+6u
I73sgqQYH6SguNm+89U9eRX8g3f4v6uUlHBQeCMloW/rT+3eGVbPpDtptkBzCYRRM75fIw0d9UKz
CUNtyd04L06guMd87yIFZSNs+AJbJHElsY09MRkhXSwGrUDhtITFuWRxqdvVpMt/7FW0Ji2H2Xth
isEvj0wS3akTrZataKqJivceelzc6qqIooeCIf77T6+SH0VpoliA5CqBPAejDlH5kBRDlZ4pPzbJ
Ntb5oIRIu2P4dWQU70HfHtQcxXJlpYJVCFRIp2oGmm7+i+GYC7XDRRBfip3J/gpiDnXAmJP0Zp2N
TIaG4AAZwa9K1gpXJQdK4F+SHycHoI9Fh+Entzr2kTPOnXqoyAiTvAyu2kWrUIRr45T5Q0FIMpw/
oXoW7806kG8AwhtAMIbpGxFkFWAqyx738qRAEiDalV4RdY8ho5XULfIRA0bs3jHSbtGOj2honEa1
coS48l+bd2kUQmpjzBoz5Y+I0zr2oPNsm0rB1EdUpuxhbaYF5kZeyRoHJa2doDzqAiJvR9SBHBbS
BhQWq+Iq3Vx4YjSyd9q107eGQQQIOKjpBdMI1zmiNp2NyeAv2U6N4+56azyeY7+nAJLXQq2Eo4Q6
ZYkxpFYsT6nkN71DFNjM3oViusmwfPysMemDNzfLH0lIRZX57W50gZSrxLugDy8ZzUUvkznEdUN+
e62bCzHZQ4LlokKn79zIW6Itc3JhdBX9yHCyfpjqDsvWQXVcmdqg6SmxEwCxxxNtQ0HL9zNv7UQY
dHQMVSgFjB03j3x7daYU/6dGqQCQ5p2wqjHnNRX5XwcQv9hoyUhuUmFUZxK6IovvSGsz2cSDoThb
aPlT141Qh0V5Hp4UFzuaH4ZIVE8yBCksnDZ43hf5rVz5kTTpkhnVPXFNo+HLLjpWE964+I+9+lsf
MDelXg4+pnxP0ZBmsCeLQ5i3cNQdW/RG8m286HQ/Q7UDV7YxQDnUbX5r6geEgjLUSJzJlXHDrbvp
YD0IFEn4oi7syFjO/roz/C460opdp4AmagErZcReUMv75tQpIx/taQvnC6aXDNy+wfIShrAKPM4I
y+xi08qRn5yJwDZ/kXvedgL2h7cEzH2YtMT/VtU0tBINPXVRvVZOeMjyDaXIpBimD65H5z6/4lLz
ABQIRqQrFOZTO7JY6wQf7+R3QqBVRSqzYpA3x+24Rcccb2R2cCjgMNbSgquazFVYfOerP1QtDzmM
IPz4/HJ8XWeA0saHVibz4bk17sMLxacOs+WBCxl8SdiY4s4Rq0d+BuHyIUB+cC8fCdMT5Isqn9uE
5Oe6XOglcMFcwsXTcCM7wHp6vMAGMDJDf7womET5wdl+64v2Q6y7JTGif+VoTRWyrs1jcXoXIlpc
DCuLgqXQ0JZfMoD2b4q90zkHpziXbYmXU+Snd5EMi2GVbtPVPLKfebVVJz+cloczQxkrPuzGVoLH
MOAXeQY2+Z8B5bVwXsn0o2GfzxzuElImBGeBlBKh9s9lJvlB3Yka5+PegFDQmL95kwLdEIqupvPI
m18eAawh99CQIrEUJS1emnUi3BTdJPw/e0MT6KOTPPJBC8mYIBs45a2vPor9cXh6aQJfbJ/U7P6J
a78Ig6Gr0Gy1Rg3rwaL+xRBzy3urRHw7TZZh10aVjCmjbWFocz/3jj8nH+g9/PRMbwx+xguVwyaY
pEwWdVAgyofPg4zaA5EfIZA4nf1V6DEeNXg/Y3qJkE2u5i4Wl/bhWh4WsNW8pUiNEH2Rtulk4dpF
fXH5+wsnHsI92gX43UK8EHB91VCIxfbFelTrcDDGwYdqGq3OXw/fZRsoLBX7MZJUvaHysGo+FHFj
uQ/c6s9hd+ZynvSGDxpm5t4/Sn9ZdsR69mE626T5eNmhlARTi0SbrvuZJS3AChZfJCabdWZYRNju
Bc6nYAXnAIxGwuJBStG1wqDW4H4GNONb95E5G+8uq5ZYSbHUSUD99BbPUgjr32D0mOhz8Fhu43wE
roLBqanjDSgAdq4e900aVULly1XJYcq3o3w/u6Yo1Xq3POs5fEvPQa62ro86odf9CsuFdiHmHxfz
gmKuoZVSc7PSzUib3ZLPOVlIJEdFlIr3hudeZ0gWe33KraFc76tBkhlX2pFR9Z/jOzCUnnyVdi9K
zS9DEtVjChj0Uv2aeV2gu1CtOYLOc74rYkx8WJ91WrkgFnW7FwYdzqX+zNfzn0Weiykyayi68e6O
PiNEyqjZ7/GK1Bam5PEVwWOQGXgir8xfQrj+GyzprvEpaTME8xFh7PhBL6mdvAE9+6dlBYJx6w/8
arD17WLOPm/WzNycYKNFal60mKfR0VAmQ6Jvh3ElmyjA84Yw3voU7npAynebEegnuA4IVS3gnNG5
VmgsB+TChzAYDTCGX0mIn36B3zOfdCx/vpFy48dk4t80zO6XtuuU4hwsyhMcXqkSwpUVnqRsa97p
Ipwpe2XtwVzTzdgn+Fmim8NCrMqaZp2l3kIUWGGZbuXe7/+IMG4Ev4l47z/Jj+UV62Q2sLdYtLtp
NQVQOpXuccXwZXN5CITTxGSTfh7Bf3O3wc/MnkyMzpnis7n4LA9fgmJ9mmPVfhrfHoWGsLHoH/PI
drXH4ArjhcraZeAJdynxwbyj/bgne7TVNLJ4GbL04K+XIlxhzWOU4RjgwuPlwKVs6vEZCKbSfVs9
oj43/Mjmq1R8lCFLGckfdVtX/pgk34WL+KxrHcqGgIhkx655XBy28JyYN+LCzSEBrqMmrakdxWlr
CC0F5/3OV/0tfHTgBNiIV4w9a9/SO1J9OlUcP/B8L9dMtHOeCbeUXokERjBQhw5FmMMfjWdmo+2r
Pnmki1BXkaI3muTUKnmUglIosM9BuF23s30ys8n8sUkj05h17PJiqIFPxBbp2TsULxgk4ltlZgdH
UOwWqhe5Tufhh0RyxwAQsxBrv88GldJpP7tYCI0/jSGfPW0quQ+IM30UgMR4pCv9N9v1JFTtkPDp
zUK8kezyBhjbjp2auzTIVVH3bJuos+m6xLUdvnCS45NYJcz2PsLuCori/P6+Cd9zNwxfm8xIHsjc
rQkemlTNUXgd8GEGXo4j9C9pEJ4seNOEnDmxiM0mqAShjZNMmF05GrABnE1oYw1UtVDpz9i9eTt4
8c6QvOvNaUeCuEg6rhkxcOirg+ZJtGtZS2DogvScJiShFCzMsGG9w/a+H/qu+KTf+A7vSD4n7Rcr
lfNRSNKMLWBEfRlKu9et6zViRuSuSQO0rntVpsKQ+Ctem1j3Pt8MZkfInKJiIZ8V216f3AyXhYTk
gLtRx+2Bn10/wtzRN2CnsMx4DOZjn+eVUz9tNr4ylmF0lc9QltN4nn5VMV2dRxtlLYIanCTZ6WcQ
twhvhQAP6GS82SPq5qB9nKMScHGeOfItw15orjFd8a0JWeBlFFInpVcRmUQqj0gRkpWRX7wBbpSK
KZxWwHzXbqhSNrpYALulHJF9feO3urDZ2MTj2EH6uoT8KkCQjMyDpXp0CDBFSykJwgTvAWp4Zl+M
A3DgqdH5K2Qkq34Oe3u5ShXU+QVyu2zChV9GwkfeuBbnNB1IOusZjfim+5pQ9w1YcOU4rv6Vv+zW
cJaMIh4MO2H8rKBKQGKhpcrQe/o4M0b8Fkfu76+W8fMmngFExQy2UjJ0FY4++kYRyo2Jdnunu4td
H0tJffnRTw7T/+0lNWjjXm//wVZvhxjbgjtRVU2V1LDs5bUlThW6INmqkRVMxy9yYaG8x3L3VriN
AViAdDvNR9T6NJdyh+HkFripFoqPGiy5HJn/QZJK8nO+xBSsuQrHy1fsLXfNtTzXWQNYUr0mOG2V
kLzco3yTodzNpr3pyJ5iK92//L5hGMBNp5Y7RewKncRE3KuFD68/i9K7cAO3ptuJ1wy4ITZ1hRem
qTL8x8AytGQ/wL6Wlyhx444Yp4w+Y/W81MlLOKUtub2bjMKkpGHqjuSmlmbjzGrIBSacxQ1Nmh+/
0jZNgBEQIEwjIJQK7l72KH6Tckq66BQs5ES7ueGyGcu53kACNqNDN2mPjhNBec/d6cJS4cNXrY9P
e1Lndin/+/dikdxfjcuLyh8GsOA5LvZYz3YyUP/dd5WewH3FbfldwTphZfWgXjRNSrJNj2ThVvP0
qIuLDc9WgaKjw8HWKvTSgfQzZy/YrBIufcLudkrBPAGlh/lCmggLoXktjWf5Dk39qmS9bfNGAS1Y
gzZtGBANCEojQifl9NUODTJBucM2RZizA+KQnL7l6CYKvCukkgKDB+vVhttqdxX+4c5TxVszLSkP
6HXuPNqxgWLdpSwpS/o6ou1DHZJGgP3Srfjiiy8ks4mjxW7NEL2sDGsA8NSK4kMjYGxqqkvHXH39
znQoQWwMMysGG069qW9GhxGdm96M5iGfHKqJGPfdGfdgpafZZpN/b9BJ+n+X8jN2HwQWwfrxHt8e
XWlYQsz8zxcc3a9czYqifKYbaMlXjkw/bU9OjiJK30t2tmRZRMQTLWf/Z3nJjJ1vecP1CPiUJCXC
GpgYHyvGvWYafKq+VF/3GcfO/IhrMJcjDFt6emOiCIvAft5rI6Ta6KiM6d4fRY/Dg/x8EEke36og
bYKjrDBOPnB6CABdveTvWJOPMsjUNpIsnq5YxYxhHhgZxBpGsOmXKQBkg1ahPsiTZ/d2zxaFam3S
elfgRPjkAOUoEYKtIGqkWl3GsBiienPsc0cN+/MG/wSupugWMAu956CHVHqoDoc5bmjzq+vV7PGY
PtNz2ha3dKTq7eNz4ajMRsuGAHnDo/+OIq34BX7b9CrOO4EtQ2MZ50fFDLbi8BrVIEn88/OgVDT1
CzadmJDvu0rImJnMWiVHE8DlbbZAw1OfkEKXKPssCvNdKBBvXKAf/zSuACO5/IrZwTtFn0TBf3s0
rp1JEr2sGpqYvb755yPv3c8I81NrZKniwKKa4//0uN9SGwofOL0Y4dzsxuXYBLc3N2kORk9AjimI
kwSI4X/3JtmzvBlu+ArDr//CaiIOiz2aYY5CQj14P7JzYD0sVEj4Ox0OGCETDVvij5r74UeM7Ouh
eth7zpGzGp/+CKwP2n+pMu8zOHRlHvd1E156+frQIh79LjArEGGAScskdd+ag81PYv/9uMb1zDq2
E1VY83G4EEkYUERjDWr9tYZh/QpMLCzApMnyuX0E+hEdBvTIjrfzsUb8oMxWOuib93tuVv8i1fQu
qAwxv7+bKB0iHo4QBWIplELNg523xOx2R5kSW62/J2sROtFWJ9QnY35rRkxYn++KsYodTv7kwIpJ
ksq3WhR0kUusjzdgVfHeogCoUetEZo+Gjq9sRSVXRDh9v2jSOlRN5VHwXVCRY/Gf2nMs3eO8Dj09
qIqh/8F/GrRLLuU7HDMpqxaSrQhd41OTAza5PBigoaFVRQynBpi6i96JXeOnHjGT2MluZ9p6az8j
DnwfGjt8mHfWuiOYuiHyNIKqb4vMlefmrmb580adLv6+Q/DHs0sBoAYVIT3GhE4DtI8ahtmUWPLm
vOUWYdfV71rDffDg1QRsYR+SHLqus3EqOfLqiV/c8zr9g/iS2YT+V6AXGfra4fjlR6B8Si/87L4c
/8fKOdH6uHOEkq020YgQiK9KPGM3gqoYQPjaG+OTY4DybiIYmbt1p2e2yE84MsOd4sMCgmmH89m4
uMHHB6q5to8WOJ1F8pafrszQoTkk/mhBzvTaUuREBOQS7HoWzLc/mHdJij+AKS9w/22HGXysQUij
StfABzVW0H7SSWhpzgs2itMR6lJmXANHgkJxJIfzuOWaXBfaOrsQ/FpeVy/8MYlafc7s6r76282a
uME7pJBt8K1TgnIfgeb/WVe6mUTPflwRL5NQrSzw5bfKCxfV2EpTiJ9mw1OLMHZsa8bGWt3uNyxW
w1avKj2p9QzQHQk6XVvA2/RRZ3GFOU/IrnHmEYYxENzskmXldqLEtLiFl6ex9WFRHguHv4OQ/tXY
He/AwhH1BZJd/cB8tD+jVdwk0NFktDnkXirVStpgkx1IFt8u8UdZ/H+hRcrDieLZ85y0/LzdjVKh
+Ksysihtaszoe2+EqGx5p8QvjnpGWuhiqegxH7866fhFXIkZ/S1jrdVfZXflcJaWNwmuIpTIoboH
Zx4EHlBrfpquUW0bShVzaH6eoAfFDsLO1iFGVIPVv1CBj2MIih6/GrEyWgegBdrv/gLw4ykyvk8f
EVHvfmh7dtZYC81W8QqKa5o9IwJZ7BMEvUIJtsD9F7YkG71+ve+8a9P6HEFZQNQEy4PqnvC+fonv
7pMor/0dE65ZWUGvrlPcWmdzfJgoShUXysPaP8Dj8Q4lctNEPRdPQdfhNLKbDBYI0muUSKW5kCq4
pMqMJr0xajaSk70Ao7CuimY+vX3jFj471Ykhwv4utFHE5fvPz/p8Oae3iEYGFmJ8bFUoruw6s8c2
iCsbbqdRtIKLfOSPGClvV6Z463DD79zlaNWcyTbUUXYrrVXtkF2uRf92aqD9tP6dyFNnKSVQJREe
Ow4SeaoZvY4fLhpo5LASO3iECXo4WvKQmb/OIa1R2RV6zd0BGLXTXnt5zAPFkK3huZKtvqy+CD1k
inUUbYEyTQDWPiH9yAtN7AaXYcWgs7rYx/qmJY0DkTo8B6sMszYQJRVwTjMO3pqFfQj0lZr7M+vh
BKik6U2P7FFDGQwNkwXZhha5KPjsNiHXa0IBQ8kDEbdA/9fwJwvxg0sCmflzKfHnScRBMVTXboJm
zehyolN7BGlDk3UjGtjPRe8I0Bb52UlueG+XnZ+rxkGA08K2px8KbjqWHZFofeJU8A1XAAJWiSIY
L+gO2LSkAn8kZQLbS+WLsWVPbY6J42EZELI1SJWahjbh6E6n8FOHE+ySTfoAr8x3z3/SOPXaFOQs
nGRWUkRkxg6pAsDEjMZ7KZsFVgzkHFkWBmtvpEDUXEr6Lx7Y2lCtsIvfZgNJLE/hs3dWtS/U5mwy
b9q1oWXZVJ/J+gUtB+kLFmE6FdV688L1y2CyPlansZYzM55SSgP2jwVS7CRNsu49erZLi5YtCzlz
ZAHoYan09I9v0iGqxGaYMhBKnagSpalDbfUpA+4LFR7Rk4PYENSheZN2VeNhr/W0Y2dqo095Z25j
E8RMeOnQMy5w/mVNvVGQHE36TMzxPZRd1URBjvjmWzxB4dSQKssTvJc8aMBFPvq4C8ldcYnq49lr
OoqXyifvBwWhT/CNCkOYRiKNLdptFT43QR+WE82maenzwXc1HcveUx/ZAJ4JMLgWTNU/VW4KfMmC
gpRovx9xhx5uJKOUvovnX+v8yciXTYGWCsemH7e3GqlhFNLpzn+JzW/yzCuLu0ElwlRJtLuRwSQX
6FiQUgR+QDGPaLseLongr2pbclFz8yv5W87vzLcDNMJyzE0rNbVxZX7LQkq9WOlUUJ5zFwKhDJXX
SAgMGWgAafQwCYDApmONCqyFLIPC2LEgr/df4lMPoWxRX+OaYQmWy7N3GB2iDJK0/1kcm7B+Lht5
m8dpB+H2/p2+xO/fDcr4cp8LwSd2ErErXrVoLpWA/EkeDroOwHytT51TSr+sALdIVzKBd++32YDi
HS6WPTqVKYcu+d0W1v80Ux9ytjMWYhOvIVKzj6FdZodEnUJMeFqVuuk7ZcApGzPwJBu4g1lpdKi7
jkPiw3N9D5ZWiFwEnfJnFLe+0A3CFESfqPOVWQUX4TBX9thUHYyMokJ8Am8sPepRp/NmWaUVXYFb
MAWU6f4zjMW7pqh29l4ATcU3GCZpi1dUAEoiBkTHsjcz4vCyokB+gZhAhACIMj+Wvyf5NFgFPQ93
DWrZVc5NPWAw6TFy8oZQ7Uq1ABtPRF+7EfKHzWepWkvTCKDexNNePpLhE2RidgNhyXlLIbrx9jEa
Nf7XAhQAtyrNLAtbIC6hmEWBE9XdgJ2CGku0S1Zkf2kofsGfPzHDoa4GshPcbRbbJZrouitZ06CX
EkgszVkGspXAiTMmJFV+JfHQqRg4CzOEMmt4fj51eJ3xyCcv4y8CXJixYFJStT/fkkr57j23b/+A
+TDjWVYvSkOyH4X/RwajtC0QT7oe3Z4Q0LA851b7awtwpqqzx3ZxyreXS0ctBlH+iSr0/YN/hP0s
4DQiEffrHYTEIF1pQD0UqkLRuxZw9h437cS5Jpa1u1Hq5YL9W+Q/aQUAVPatolz4sj225QpDODdr
CLcyjr26LAwORLEGRoXYutaYouaddCSatuBgVOIjyaHyq5IhQllVT36lRZsLwdqWh8yxmyAQFaAs
1W9FFNgj/VX+5Cl8/B3zZ4u4p0kWOu+4FIMwrxVQqtXTRzGxjGBLaKZEwzIe+FYJAmAVe79AiNAY
nKUr8Z1mN/pBHkucVhQL5XJ+5u2liwrt8tPALFMEpSiefekwmAx0BWFNuVQ+ReM+rR7vc5h53xuC
IPxyEDe1nVPkSfbdYtuRTWhZtrSsX3DLjgVKR3/ndJClgzm+sN0APiPzNHrNu4Knk1rQcztSbwUM
SL88TTIU3L98JVAlF8sKkj8x2HSuXKQ7Yhd1UwJSkf1CNg9eoN5bY+k+3/2zTsYCOvmkKdsmR08/
GbE5hPxVtJhcr2+F/yxYTgYPCcA1d/eaR+GH58DSKWPyjWrqLLOWrQ9qj9PUBiN1QFXdGAVUze4h
kRtUD/cOFr4ZuEHUk86TUTp+BWGglBKKYvcxGPwaUMdqXcDUM+yXAx93RCorbDidnVP+x2jicmw5
AqDn+6lY+S8ISPcaijWyMBYB9JcyvJpcmi4unoi/vAbmeXX5MphQLWUscwn3iUnxCjD47wm863tL
k7OJg6den4atjINReK3OIBnmq+bJfOQix8UeHPirwfFzuFITxVPZSNlw9BY/kJRt08Zr9Kb1ZCDH
3gYtBSmIdVnctSLV6wTTRRtvohGnYMl7sjxSaNku8UhHSefWolf5EfeQyi9y9RqCKA9pliR7WF8Z
b05unPz0PKLgmZEAqa3Kz3gyC6Q7KXMEMRLxbxbTSxXJ/ySDqeHwrOiOFgD1r5bluyx8K2xHiNEQ
DahFiE0hbK3FQ9BhYbRuRK7RF/VK9+WNJ1CWBu8R/s6xYSWE/LcTAH7NeCjhu76BmHnDqXMiAYhN
f5D+zEVJ4jdnQ3MPExz0upnSCXBEdHkQ1ZBPt4iTIzCW5i8H23RdLRJm8Hsbo1gJvlIS7ccWET2J
/5XY0aVCzmPpaIIGUlOa7YZgujNcoSOhvmnvbiI5LC8wpde/nGR55WaJkASP2Dv5LHklVACXra2g
Cs2t2kQixCWIMwshbsY4THbzha8PbUi0Q0pVEaSVrAPYRnLVBaV6QQ15mA52ww/wlEHilN8Mq+zT
HTMR3pfQVtUtqnaQpGEznnZsQqksI5wxyn/iiTbDNjdG+oJZVQZ4y4wp+H2TI1T4vf/Cdt7lJ9x7
aCHl9kJyd9i+jLVlTKEqTzMiteOMrw6qTYzGTcsu1mXnYAnvxME3GmP6aVKF1RGsQOxBcECsmf9k
C6T5KeKmp3OVa44tFDOv/Yf8ZlVrvrjQmuJsbHjM8+8W0mvRB2Hw5CI60X9y5bv2d+M7m8DGFa4N
O+HmJgMiug296ZRsVdWKqSM/sGkRyU4lYFn3fY3Im8psOMvRo/Kmiku2DnwHsN6WF7qnuRkM1xZa
xUCC8xOda1Z8sScfxs7hQRr56rLMixh0q4V25LEYhHwxbGvxeiIo3fOT/7T3pXcDWNY5DnnnSHcQ
HyuO3EhkWTe3PZudzumqx/Qa3u47HED1Ar8HDL7BKt+XlbEHUnZo+3l8yZ47ZxZ7OuuSIx1V8we8
r0RP6rERhj0EoRSgptjGtHAPAISPONFKjWslO39OHxw19A/9nbQqq2V7Q3xFIT8UY3XwovYpuZ6W
7G7X2oN7y7Rix5xgLKQW5f7/tRsSRAbK7TU3fnqouCGUVgIS/6qI/+NJbTp8Fh545o337ll3SI/4
Cnw7J7G2SojB0EwFW0gQh09slEZ6RBaO/393ErYIB8ptnJLT09GJ9prX1boIHiAwfWs5JCa41yWr
Sk/MI4hbyNZrwv4cha+oBmyM/mQVX491pT3tko4Uw4XFhUwo45k0yhDei7modReGPmBaQQugKJr8
spUULwvuCoa+pF5ZVBcxwkLc87oO6W8G9wFZ+tA4kmqo5zH3kgzRLALLWzRqmHUGEWkr7Z0Zqd26
HPACfswSf/OU0wpJdfRyXcVnR8/Vh7YelWxh1Y7ebVSZ2Pp4J74Uww4t5KLYuZtUTqPvycvMrhEp
z07uKVs6olj7skCm//7mNuE5TFRkBW3bknNKuLb5gSRbU8nbjNbMB1kRaYF69BXlu6FuuP3aDlb9
1sabQqcx30D4R+uygO/2hX/erea0MKrXa7YDmsO0zWckgxXhG6m+ngyE2w2wAwZ6JLbn+kIUX+TW
GdgnsUMxf9ahNHHIyvo1+VcgJUndVDMYr7cTrHNsM7C6fVHkmM4rp0mKpGvL5JfoNRuQ1dZjHwOC
OhZrmvla0JWlfIjN0UReQCyds3bU+AwiDaRWga6/nExGP9BSrA2E3G9A75hKg//aDTsjOIJEjLkr
yTvRFCGnUds47zqiH2DlzpdAdRfv1H8pjySL5mPUqOGdPKLz86vnKwP1ww4ah4JbG2hUmtnRprfJ
dRdBVUPvBxUiNQhnebCXcYjQap4gV9RFk6r1hD3+JQr0ZSfKgcKKuPxUJTmeJAZHGu/EiFVxDHCz
164T868BhvyVtSqKRx52ZnK/4LRWq1ydvZrieuggY/qzhY6F7O78fVRIZ84xw34mZl8fTon8Ob75
AjtQbOWmHFMh40SMjL3vZZ+hUQnLdx8XP3UCsj1C1IVVVXVjb9p5ci4S6myPJcFisUdxuKoTeVgu
brd4tXHy4twOnK9fpXqpxoFvdFU/vRflCJURm4GX4qbZE1ZVPOmQHxJdWKdhm4INDfgTro08tY8g
XLm4sbW4hnsjVduydMg1lqymRw8RjPDTcuNXN08gKvTatx6TaiDGWFZ+Nkkajsgj1hkC/yLXhAWT
1y6aevNMiPZyY6mm8v6hxqeZQQCbWm/my1xxQjJbzVIHe7V690ntuwAIPkQ1/n1Ma+ycm4mZBLdV
grpT0D168FfF5GEnbwRPTHSf4zXrYc/gxBA1uSgvdgCJJ+yshXSKyP3upkfIhDBUHCdnLpBtk2ne
pAoYX5nz6Y3uV3TjXNy9tYpeeJb68XS+UUqheUlltLD3l5IAjAva8Mt6mKJvfREgWK/g9s7OuEFo
tSWfrJgEORWttQIduodVAk/sxamFpBOKXXapaM4gY7Csu7oDi+tUVF8IVoqAzkGF9whLsBjOi4mv
9/UoHh+/XWELRYw/34yvZLFQpp7r1ss/EP8R1RLC5fSLBDZA1Mmpx9UuqUht8GCAzE1hTAd0mB65
2qurgZKUIyR20k5Xw0caByjRgSXeH+hebZr0PLph9M/jC24EcV/s6lf8adbSY6FAfQfWXfBhzsax
VPy2yPi559KU/cLuzEk31qfuJGviz6XFFfIY24c/BNQ95zVYyF5Emd/OEgVYtm5DcDL/wnx8kLYt
qRhO2sPlj40Qv8pB0nJDQdGj4x8HwHwO9lwh/cMM50q44s7SANrXcRZRZHHWsuzkFQzq5MXtgyPc
7lswwaT4OTtUgP0xKlCqjlXgCD49Wb7ntFlZFeDYaPS1q19i8q4i0ExuI4TeHwAFCJzt+wosGNJH
jzs71oP/NuiFpqQed5g0VPpqXZtheBrut12d9RubhRuCwvmx97LOxFrFiZ46/qOdxk/0xiDZw0BX
nNS/jfWtDo9I+EOQUBFgR49KM7zmJGbAmeciJdifdS16FkBa52Ji9NMDoFE4IP4+GA6/WoaOhBhB
5dA6jryENQG1AWUo1Di9DePLX2/4kNbYZIAe2JOAdY4/F2OvHIQJUQxwY0NkwfUcSl653TPEwQHY
Lzb4HAGk/jOwQQzfP6HYXhBYgP0h7KL0X+3E7+f8relrjD/RMWO7dskblYZo5BUeqYXtZ1JImu4P
jXeOiqPeVTnpLoRRR91eZENMI5EaksUBcl1Bep0paLWGyktnjJ65BaA9buzV9QDFHZiwfeIJMh+F
ySG4O+f00JMitTS1I4bpSAc6iVNQeSsYMHc8x+9jr1+Xtg7sfIyO6ecNCRSYHUszW7ivhreqGoYO
/PKc4oAMZf4i8pg1HC9WuHN/Rfb5cMtzlaO9n2fph381wqHyInyzToZpfR9tH9uOed4/nZUVv/44
4cRUs+qnVaDxKxrQpE76OoujaBccsm5vmMEvdlXPKl95ygK4prI/agKOcVK5YaflqJ4BgAQ1Wgih
b2qF2a+m51dAM9rAqYafNaWnx1BiBFOJToM1kRJdLtsfOzu1vKg7l/1UcJ7i6MEbNNBV45UzNPoR
OgoADtnaF+Qk20gjxlrMWrxLkSwlfgyQSnVXO+BQBYvTjOGSlcS3TZ3ceMvNG+acY21Z/bw7ObsF
Fqdvs0H/o3DBhOoT6LP/vN8VE0sjWc4WosvNVDvaEl+1FZEq7WyZ3NGVoY8lVW/fD9iuPMs2dTyF
G9Tjazu4KFIrbJnZ5TtCQXcEkdPguUMbBPBv8MM3YSTCYSMFcgXTP9YR/ZTw3TU/7emWAXSC3nbV
hZmoyPdDP4HYWgp+oFtIA/Fjoh3mx4PuH5uhoh9ShfIlrVFit61yCOw0dL4jtD6FdLcr586CqDCP
vJrsIaMOAL5hrupRuNP+kMWw916tVpI9yHMdxL84MM6feJZm2aonFuI4QqsU/0A2kk1/+ySPwTFP
eOUlrVEYaKM1GaDn0wpAVWafFzCajcyTfmr+B48wVQDujrmgLE+E6JGv5W9RP/FXjHw+J2ovLV7X
hC3YnPfM0DTs718QqgeTvh8lYHflUZSfRBd7IxTL+KuRkkV1gu0O2THa9O1YUS03g5LFzi8RnEFn
vvdpMjHKpF91yDstRNvNJgTYWV2Fuz0ckgMjpI3zWZoCiW1OTcHCFF8Na4kAYwWFLOpIq49HgTOb
S/nLW+yqWQKTDisxYRkz+Gc2n9445gftCZccwSwAAJwEsdrm9DmZRNSUucoKeTi+i++tlXrzLIMB
wXxOl8r5f5iEMfKGBY2kpOXTtMSz+pDohSCW8IJYQkYM2g6lardyvw4S6ULt5wl0Wqt93ZP9YdT6
qQZ29KAEqVHyo+3W7K5x+CAiY9r/qB5eZm6nU48yCbqNW8o8qwNOOu0rD6vzeCyPZKuAIc8q4aPn
5go4/q280lATlF43+1hAqdStDdHWZleJon4I3YVYDl+BzxVobq6OVSvrfR4gbU8MX4VwfjxGqM82
XarwRx5Td0xUbmol2DIUHzjDzI9xEsJz7+6NRwlqU1UepB6hX7DLxsBvmbPZIumCElrpFbUQLd+K
oy6A0uvGbv8sGFPWbzOmQmaT1qigzqOCXbe1eY3PaQKghdqvcbV3LxADGNew8HaQNQG3hOOSLhkE
C7A8HljFlOjt2jHBEhMRfgrtL2dplcxiZVdqpSWgziOjpY6mcHCAXl6Dl+QzREB69jnKL+ZGZY4d
IpMJzt20VXpE9JF8OncgM9mxeRyXhbMYwjOKVVtDsjWD5VdOuVlVJP8aHynjNsHnu/wK9C/39ZoB
XKYq3KpWIsV/Lj0EU2tHelIVlm0IH+TR1qSytgOssFiRON9NYNzm8yvZ6G7v0W4aA2Q7Up5oFy2x
1XiINxNkeFQqMtAs9qRbX4uQEfTrV7B2EshdtZ+qNwpfrMN/L2AN0bRj/olZ6pfFSoQfeoqFIgEX
Vf1GccrPTXZPjZTdOIDfQxRRV0Ytr7yzw8Ae5aeNjgSVejJVpihXcIpmGGib7RavKwVjGVyYu2B3
THkz/iMhK5AQhxrc5fDYMap1diR/RXMl4F0hnOi2oQfKaWtvsDVVxiPyx3D2cS0ocDFLrOs7c1db
/oRb2vVWVr6cASdhkrgf/2ccHKvP7bT2HaJj9Ozv/QNfYwm+scRGJ0cboEVYTD7mHnI9KYygmxGh
/iaS/PQwBHdwy++cH9/QNn2Mlb25Wn6zC7q6FiVE4jR8MTpkkL5MgfOoHogiEeuqq6sPhe0kFTDn
UtAci/0Y7/NIig/IVC+wdqpBob0IzAfLce7LeM2K97Z08lED0HwIvcofMTIU/qysO5ltdEMdKagR
QCkKOPSQDxsYPA6BUJNoMoq2M4D7CZ7O00soEhKcdA4EbWvQsk7jjonVJOa0oGSU1XN/12LGVLLd
8vX5alt2tUzyvu6Q0nKBaH5PwyX6FSIs46qF4INXGcxHeg1Q92ljyxmyWOSP9rDuzR0gqu8KZkfD
PBSbIvUHwaJygiL6l8mVDQRORg3mUvz+qsQA20w19eFw6nAg9/Vpq/YZpk8RR4UHkUnnH3fpdcbR
g0j1Ls4zZOBkt8WpV+7HyN+DpsAqT4613sC/vB0V2ejAnDPyQiv82ZW53heGWYj8MWulEIslhsnS
8fofYIqtTPQKz2VU0oM8Fyv16XMoZ9pvjLD3qr13D3OzFYlSl39lFqsPNFoAVLY/oRY0gDmwVIpD
bmw/raP0GpPFHithjVgRLJydtSoEYlsqEMeJQky3a5pjzSJ42QloTnb/3S4GpE++amD5tcWbV4zd
KYaFApKLQR0LgTPyBOEsKfH/gVedgViXjL1alRJxi1SQ9KhMxj2U6G8XsNCUg0joqWkvYoMxN1Sh
hJeyeNjD/7nCudNI9bglQ43R0O98YA62WwzcYJCoDpjQ2t1ObI1oDwR542isB01cfsodo/kDuC0W
fI5oNjd+GI6fTUjlyphLAJay1CzghXHLDjRsOdhNBdUvGu1plWmUj4LKHy8rWx2Dz8RGTtaKKp0w
LmUeMtV20H9LHlajOWqgmHIOZy/+ButwZLRlHaFS537IwzIL4Vy5llxEOFRKHM+sU0KIw7b045UJ
Ve+ANCOmeLafbT5cfrLHyMKdWLX6wzLOhpxg8+4etlShjQZ9P6vsEWBGtUOuN5je0lJaTwgvXg8D
/3aJdDbJ7RDXJepx0qhx1gQIkVHVam2QsB5zLFMWNbdYWlifv2I6eXazMrO0mE4b4K/dyl+cpWXy
rfPd+4XjX/HWY7YNjUEeJSJJdnXLZ7myF1krcgmbiGJ2pF8pXKxEIb9HqcGv4MSaV8c1lNMGwWiJ
Awr1P6iDprIp41SljSIjoNdRwX/Or+bUK8HVYZTKAPtdN37jRb+TLjIh5xUMtEjp9DQoLzRniI6S
vOpQi1QxarcERcBVkgjhavPzfznvhXvaOJYJAC3JeicCUy2TSmwUkx1Hcls5Ny/d4XpRbzv/CQQs
IPvqVv/5+J3sb9EULK8BUH54aspnwJhUTD/onDLE53QNCX0IXeUGV5Pz2RwnvTO+zgQDHUvUabIO
SP1NzjSg8ehV6upP/el6Q7gAnwbqxPwlNCymHH8GG1qS3QnQXhrW09hnuMr/EvUcw0LB7Fm3GGbP
7ZHwYZACTYQlD/7cf2TF47kcJC0QVe8ireOL8prwoE3o1++qY9tsp7w8P19kUuGAZzC7cH3UHVK0
wosj2vpJNkni9lJpZ774sdOv27rU2qmj6KzBuZCi86BcKbBXPccCSHl+pnUc/Utwx1UJHPNYFWdo
9KlV211YX+2x+0wO68I3pB7tdgmZh/3VWDKv6OfnIgeFk1raBpvM2pi9XCrhymh7KhGp9hzbM1QG
WCg5iJGwsDLwyeoJMAr538N/oaTc7QOD4IrAKin/nNMh39hc9+lUWpjoFWmUBSA6UOG6FCfUz9BU
+3dGAY8ShQ4gyZSy5e+7vq8r6na5VLBAIzgtmHla6e4C9EEM1u5bSMnS66Vy612jRhHhRU6gdjlf
8CvFjwJPN9JeLx/pM0fmR1negBxfdIZCrRZP+3Lj46wbd1433YIhhNa/t+FMciVrNyjP4OGYG16/
16d+b3kTSJ6xb+jbLWsOFH4a+wDechNOlc2GkauXJRXxNxJoDC3ixb0CafLQvDkwMb9nkmH7wh4C
qh4l52KUB/AUlmK2paUwT8pXRH90rXls/yPZwZu841gp4M01uYi5PsM85NqoHR+uaKN99uwnhWli
CD4i1uxQHKQSo3wD1r+0YcqI3z9IIyYr03Bam0I5gIMPg8pJYmgQshqPaylvRCfn8PtjAACIQ59P
VfRFmfoELgAE5nKH9GRl+cAcOhQQgoiDQj680kBCQP0KIqOhi+r0qQ5jD5UmnqlQcyVJnJO9XU7H
6hQugJ2aNugLdN1Sfk5Pnu8M0GbeQB9Ie3D+0CsX4l4ogDNoneCyWIZWc35a3PGd82axOpHVUXqr
46uPwoh0FfKH00aYnmnpJu36fKwDkDU57PJwEFDwbpKqir71O0tzXai4IHcqore9E38SYRz45ySD
K2MZOGrtOXaWVABZk/vzjnNnzvx+zcDipIy0pWL6mTWsc3XDkPj2w4AsX+TLNZeTvdXPnCHWA7R/
llegBpoim6Cqz3EcGSQhRPdHK8igj1KkSaVCIFyM2M4inTzopb+N64/OZYXnK+U3ii8yT2QQQPwk
zVXW1iwfliVvelhVou0OU6K1wfZLh/x/TLqgr/sxcna829jkX9BUkl5VoowxhFali4tvFLwm/TAz
7BYC0NY4K6j9i/UEulRpYeqsyysSgnpJdOtelFmw4Y3SFJv83O7PXNTvnImypWSA6X/X06V8A3Bf
ZvmU9JSF7CbUg8Ib1j8jFflzNGS3HqKWjeznKjlQjsBiJ3uS5K+m2+7u5cY4N9HeukMdd6WDZvnV
PGNSKCaF6Wd95yVbIzJpHTzlTiD5p5hC2ImIYoi9pJebuxSHDPn682YfBAOZg0sLXM7TvQIu7d6+
XSywMxQzaQkN/3HU1/9MeiHlLRaY+IKmZEdnhGaOpaLB8nIiG2mVbDoCODcTKen3QYFMj7K3ED4L
JBSNT4qw0zcJNJC7eD3PZrJc/IopiFVRyjf8UZG/urnpPkK2pH9/d2taI5l+P42hCkH1PxrauWZK
uAyVedpm9JubOtKfTp/LyOFE81jXLqWvq0TKcWpmC+DyhZLtMuErhzLaLpEK4QdNAo81ghkYySt2
jflPcRscsJvumnfhClnggDg+SC6FEbbV6Uuo6QW3YRTTb3fZwSZFhkszN5KIlvK/f89k2+9KY9lw
FFVvJYCq77QdtWwLz42pUK3JyQdoo+vZ94GTyjLehoNR6+7FL/MIrsJP7oL7LScmwRxjgNGRi2PW
QopqqXileEOY/IIXad2cUF2VUagMd/0MKr4U8iZDmbphCNZQ+02klGmSfYWjI2QoG+tenERKzRL5
05wAyQkVVuLZtTyjxdy4rlDh6iM2Nw2O6j9VhKIVfMtq0YrxC7s5SAdmXHLdysyZXaqBplDPbciK
Pl9lRlxiHzpWUMAAiy2ioQ6+SmTCffZkwkrmi24UcxpUGln5W4vd66NN3Fb9vFYjSU0WrNKO7lGL
jxtdhz26FSEvtpq3rJ+zO1DjIG/5l2j3mCU3hGep5MREu8qPHZ37I6FM/QrysP/0D2dSU7txcX9k
MLKFCu+BKO82k8E9Ah5nWtgN7oM6vlDWGcXzr9u0ZmW8tDJjNGsfxiG/E3/zBB22QcP1BNUSnQ7i
yR7FAuCNtFgb1fh2S2JMnjb4MxjsoTsyz4vsQoKG6lZMx8wzYBH1pNrtOXQWssaxZhRAuxB5cMJF
hy7W/EH21WgUIpI6Dz7H/+AeVBrmuV+bSlvtGGIJBkcTlHFtAvCzBo1SYbd0+asK0eP7sUK1jRAK
Za3dJNvTmWY1i+zMcmMRkvGHG1NI4/dlcvI/6qobrQIq9DTyU2xZQw9yUkuxapzx62ePjxU/jdtx
S6RIGzSQ8JNMReWXX4cEc4+0pz/Dt4hLxk9dplGRLBOmpnCSk0NeFX1htQyHIxz6hFvFAA1baDKk
d3gEpivYEhv0YsFMhmQdy4pOpI5mnFUCIeupky2gOPWjOX+pABFB2DpyoboN+9VGo19ECXjtC5MB
ZbTQIMfYrb9nG/aHp0XuzumoqUk31/wiyr+ob2dLIjrnRzwLVHvp+3vkhMcM9QoQEFpT7Kzft31X
b7FhUnZVOb4ecgIfULDkxs+dv1zj84BGSiKklvL0nNeWfAoCtNl6n674dEMyU5zyl0I604qrsj5Q
nzy3mLcIwbtlLVSxyckISbmJdCKRnloKMm18Ydq4lDEJc+fMSLHwcLjki79nttAfhcs8dKDEJHGj
J6WOl4vCee9Hab6WKwatAfSx/ZeB0CzMbmoRfAyeERNI3uFkkunFi9G95aFJKImQ3IsK9TQoZiJ/
8o1G3GEPfqCs7j3jOF8JIpLtWpGDSjeDlgNB+8Hn/OqwwgDvgu6C6QMdv/HadQ84RFldiV4HaP1S
ByAVYJMND8CEdmRsygM2XgErxR7lBc8E51UT6yw3/umeUY7uErYgkqk5hKi0dTeCVCtoZx27EKbe
N20/jWb5yjzIdTkho4rvNfme4Taz/Twz1ENiomavf6ohL6FH7rRHeSeYnL0BUhzSx9TWzTPXUTFf
wiSmE6Rw/7pqG6A2bsGI9VkNgAKEEJCwNbH5mHzmYE90xgzt+jX7OHpgKVD4usIwpNra57Wg7wKx
aDb5V7UDBRAx851s/O8QWp0jK+rRaB9MuMAOoKKvd3TwGpLsZC+ahXceO/DLV+9PVfPra8mbvTOD
xb7ppdf2ZJhEuWlYl6moSX3vG0sDLax6fzACxvEr85OkXa540MvkurH0djU6qbZeLGt/hoIrU1dF
O8N96gFxILSKRz9i029Dot0Ewob5IVSuYtD2tq3zdjo/fQtFYo6SThAFhYRtZUmuOEeFR+TA0KOB
KpeHiR5g4zwXRpn0xq4mxqXoNrkfP+6px1JZahpytCXVWZGSWtrt4NK8nCtsq9OwRfBk9Bqo+3bS
6C4LdbbzXVvnhj/VgVFPnpBzOIpJRdOl8bjgvXQwn9KvwfWKVR17Hj1ofyHbhAqe0zlRtPUfVZwH
/1DbOBXj//4p0j/fqgXgfCVimwbjsFDu2FN/7+hlEtqKZVxVAahUeTiW5/GucZ2QlRq5n5f/PIgQ
yIa5fV4+2Bjj1tWCg7cFKWUb1wDXNgc/tNs0b+o7bzJ8HROkCDgkCli8Lj5VinS8ccltMVTauXef
57xNdVWUbso68hfu1I3AkQb8m11ScknujXZ3EfmIVmP+iN8ZYjbq+Pa9ukNcHkz29hxAtBh/qNHN
fmF6CJyADoGN8fWmLpdpysyffsbvFG1R1SofREEmjLjzuqwqPluiEEDZ9uHzGOwy5/CD2VqdufbG
bRnBzURo/HpJ9HkelClUaQvXl54ylFLN9uFUQjuqY1aXbJUXcBCS7dt/6mr/20it8wFttpR+SCjh
W9h94LbkbYxAWzA6hBE7L4IB6hhWklwBd8F2UwNkE2OSjyNRHrhqy+wdl0cknVbK63rTbmpvmNfN
UtCR61nDbrlIvJs6Q7NtRDEZb1BGOibPN853d9FLArKqgndUsh2f+JbsFTfWn4/xPYz04Upr3jd9
yrszyzkme37ClIajX/hc9XVnXEavlPQpSif5Ff3W5Q8y1mA2YZdrBdR3ONF776yhdATsbg09LRdo
Wf8/soEWoQ5rR6/ds7ApjWYNi+ACUVTkAjbAt3cXmq2sM3+ohHivDb4V56ppkzWP7fftiQJOzUvl
ORW1RgoEdSCJbfiXryYYWlQHhWUDXtu7FtlgN3KS9MvDGoNmRBNH+m7bd0ndtShlH2t+tDEBPXZR
rvMab+GRk/8bAvuIpub6QUkqrCGKCYuKPMyGUCtchFgj0lO+TRKol75AUx6ZJtbCSGaSnhvjxXEF
e6c0ugnHD+YfsQO52F700HCNr6WKuIPUq5A6pvCXFH/JoMmFu5nVQ8HVcAZElNRVFq5fZOY5KCYy
xLn/GZTfpp1D6bfn9r/mJiFuQg4ydvRRZXmDKheYTTzzYpDH8Wfh2K5buNo0LGC2EdveaQEbBamy
qaPG09F8udInBWmaa01lZctVve7irFd3Eww9iWYxqOoYyni1/QXmDjFJF2yhfX8Ko9f0Rl9yydxY
RT6rhkPVeH77Q6z8SXMSoCE1kvitSyFngY2pFQlh4PQNyjAIEWd2U1uxgFlb/Tr3R8AFcRs+UOZa
gDJV/sCQp+QqptZrh/yGFgwb3Vrj2G5MhzBADP/FPUXEjoA/22HOHgttiq//Yc69Hs/n+92pTzgi
gH4af1mEZyCArPFlgy8W05VsfcT+gBOY9pdbTaLUPRSfMz+T3A7xqmeDePRbUyT2W6/Qv5H6c6ne
5TMAYujZDZKpAFwoJhqhrxN+YfBz+uEmB0rcJ58CK4yN15m+wQzy85Hpb1kJ4cGUC83jg2YBF2cs
Y5UjXCb5sDrEqK+GPTVuxZbKjgIvXbwlU2V3wAgGrwZ1GngwNChum7HVtu2mg3r/qrmksOGGNrQq
pBvHkBYaQUIUpk8z5I37KynCsb+Gy1/YdjtdIBwFkatUuicVJ/2EBnUzDIa0Cs3Eaa6P4hWxGvfD
gbXDFGrsvXxOz+Xv0A12q+cY+KMceye+BfUCQ5c4oP+vwT5ghgYt4i3zBH9fr26CmN9kIkVI3nZE
faa6jQjqdaLREP3eMWJIgRdAyBx5OgbNpgwAAanYiHXyePNfuE1ZXJcyZ0/yJdizn8lOF2uEz3Dw
0c14UkU271IDyXcv/hoG2kzGfUv/4SkM9mqIZJnmY84jCfDGBqh17fYhlZaUDgyq8ZwJ6Wj9P78G
hgPr+PNqf3yFG6FxaKxHZBFdxmH73o29DMZarMAVp2gdt8WAggl4Zh/XKsGKT1LpfQkhYYyTZqc3
8VbqN9+0qxiQLPloSABTOf5Z19lVEvlF52s1vYhDe5gO505XxWsd1HKiyaRMonwGyzfG/6RoQH2M
Y6xy+MyXTnAhhFNtar8HA/zMf31zVip1ISg/DFmRjtuUPkxJ+tWCffo7QCP7mftf/tlAnqV/GTld
JOVpmfz/U/LCCcD20bZQ/9SE7rfcoHa0AqHHwWlwQlqAlKJS08+bzfRcjPk6m4Z2nalhfJlE1TEF
14pLNVj8xhegGRA4x4eLezJaZNMi9x+6/efwjU7HeER/HlfPRDs8BXg0BeLzhFY/S7m5fL+k/lXe
+KKM5rXm/73JMu3a7Wxgc42gpS1pEo1gytweOOA5jqpTNliJ4Ss3qQKu8neWNE1GxWZeei9dtkP3
CPortO3copltHnYSccUGbGcbExOerUv19sUzfA8GzWC56L80GVpaAwrw7227yfs4SDk8CBJTSOsb
gd6yTZSTYOwvyvPhw5leM3DSzxz6NNv7DqLwFfepOmM0KwM3z7gPNKMbV0IyU1A6EuWacoMpl/0q
xhn29S+UdMJ5leGMVY5PECH1p7J3fLPLcuzSLbo7pVSUs26X99983r1/DmReq4ev+LnGXJHJpGCg
1kNQtJa+D0oThwgv962nS4g6uX4dR+aS8J6eLLER0trJBzqPPkwOe+5PsVT5n3rtV05r0akvpNPV
8u3+v6g2AYimVrtqiUjaz9py/FqS2YpXCpscIIGvIdjdxWwO7/5JFjaweicuu2IkzEeTdP5duoYA
TXEP81FQ/tEm3JGg9ZusQ3H82APLPIZr6HCmnV24SUbWgkiLDvxrJUxIs3OcSzRv0kgFZ4Sem2qj
/5isAUQOpw6qOWBoT/mW/UdfhsSIPw63jAWcC3yTXu/voah8Y0PvkRvcwT4iC8v5KRfygklKLl9y
a+5CLC+eh+UOXOOJgPypZOgAIvIcJ7C7Ka55du0+x7+9P6JZ9RaH+WcsjhCbfmK4O7GbI2dXPpUw
YjUZRQy2lpSvYq6AQLcFCAA7Q3nofsCG4rDY/TGbyR345dC4buQ4T9MFO+9nvRxsywpZ4Qi50lUM
Rg+kJxhyJdb6wrSZuPaSPWx1gAoxiulUx9oxMhzrWP/n7rXeEuRxMxzfzk27gPhs6/uTuxuC3UvM
McGbs77wxRyUaTVRAkpQrefpPPM6CgwP+jFHN2DGEDesVlOogW9ZacbcZ64jTd3CoRIkZwwdg4x7
V7icpnWGIIJqhkGqWB2qOw6K6xcbxeqBxqHwe8gbqaDGNkVS/lzvz4NP3cnl/VN3/xaIAMVENOHH
vrIjbb8r6W0SIXrV2x3wx2OEzVGfKPbW75nttQb39+yP/80/vtqsN5TFhvaQx10tjrVQFQPKpGRm
dLl6js/QqJ3pmSvHV6DLxHsPK7T6pkQkf6NkiySo0wU7XMw4Fl8RXPbDQPXRLngs+mYObuyXL0SE
nC5KjyYmmYUkXLrHfWDPz9XgmOmy4WbAWH22u4CNlCqCbL88nM0ZGuUls5IzVx1OE8caDTZn6XyZ
fGrg0CegdnKDld+iCvGorPZtvT9ghayTfrXytGZX5FU6HMMWRqbcnEW89ez1Hd24ewZ20X/I03M3
y7B0VLysBVL1WHjUwlBcWjsx2oyNVYIpOiUqdzVO3uMg6qx9iuYven0KrQIiVY4c1943F4NPEaVn
6iCouWH+7iB5FVCSiqioypsEL9zEFg3doQqTbdOLSZa0J4NJrs0cM96DqMjXsrlK2Z1KRxAorahD
lI3quowREU5DnDcZtrtSaD0Sd8/LWRWK87QI4gBJ4zfMfXjyKyToxGXcevePQvrSrgZpyj0qTjsz
8yrhPQUDy6W5HVTmCulA4HnpP6+blR+ttJrlBJOJBxHNscuqQS9iGx+HjlrzNA/aSJ6SQCx74lrL
tzR45oyvPHcCs8jk6Wn6M/3GwxktX+Buk1Z2bAaSqd0i4wjffwkh2SEiExVSWSQOI9nLJqapSIdd
0yUL4/X8Q8pdSYAwRn3nRfSdcXgauRj/6/6MdmyozKBwAwdvntEHKa7qYYhR4AcKnqVyD0KjjlgJ
bgdtakIQ/Ji6jRSH6ZXu5M5Tuf5c1nPfCP5c9VRgWZRGu1fqncmuBj5ZtFR06QfmizjjxLKQnzkO
tRJQ00pERA1aO/7GsKZj9/ySDJkxqtcWqTBE5MU+mXiMkOPwzJFSDyuqxQRqBb5f8Ofxm2zA3Aip
/WGipYLM4Kb6D0YPdEU4F5a9OQC8KwdkP4ezOqNuzsE9Te1y0oqxlaQgZhOhDwyA4ItBNFlMJbOu
yRptoHDHJC1xJ+KGKBjakIAT6WmhI2DBn1MF/ollW84T7Km7CRjRthLNgjQVzPuW44nJgE7IW/zh
OAuDvvQ1DJYqckEBKIvwrhDI2HVIpMa4p9QZz2our8fjCr5RV0qTV+eS23jJ1pUaIpqzdf9xWMfe
trIaL0wxArfsdyIYJV0mBXJCsnTQ5BnZNHY3VX6z2rXjK+u7N/ICu9bHYvp+SpulRSG6+RLbCdIp
VIEc578/X6R0YFDnO9t7lbFPaXMMDPvRhhrKmLZXgJ0XFlyrOTkCiSnGs/l1i5jtQ0Mar6pzXAWT
QwqBHmElEj/APr07XuhqF7tkUX5RTDdK0LzQfF18v6qxBKRfqUk4BeEF4V9klqKKXRjI1mMcgeZT
RZNBQJoUQO8xRuWq1opDePNzUxwp+YGjCwKWHY/i30FjbkNWHtCBYcAIHn+L5/GXcOOicL0fRRji
YzXSQm66KhpUceClvt0dURtrxDu061shlPoQ0DfETesinqcJ/Np2wfKOveFmZfpbcKBCARRTIwwb
HYGrZQx7x2kfgfk4+MOMbYmH2IRomDH/l3N7TPX9klT+NWTVXvU15NCPALOzGDOcfX0Jr+IEkrWb
0igVZcZtdmOJ0yZfeg9d7aL3XlSQKkPWP2FLXoWxwgScFR2VD8ZHtcGRzaAwBWvEaNwm/xG5nfoo
fhZ2ugjnw4GULcwLdgEdcCZR+w3wXZS0+EH+fBc6hqCTPGddBIBeQKEfQVTq/X7OVB7J9Ah/RtDV
24+VQ5l6szS7ojh7nM6ieox4qEf/+oi4vKw33tMZT6UDZrj6G6dcJqzGk4JCdSPwmlYhGDUd30Zo
TR9zMvw0T2i0EV6cJdZgZEB0I5o3gef6KMD3lBynoVaLiW9fwZCcflmjLv7CDsBjB7x9spYmcyQ4
B6SjWO+l/TQdPvfDKveoSOxXTP/Msh0KMf8RVvA1GXB49cI5uKQzR1p3IMh+WSgmQ9z2w7ci6lhq
W6JN2dTOzilB0enuTKmoBCaH6eU2/QD1lryC2tenev9MiA71mNXU8Zu4WEq4bVTZlKElbU5/69W8
JJSEC9rOmUQKB31RQ8El/t6M2AMPS49nqoidQ2+yQeB+XN9TlPy0KHRiYkOg5Cr8g7bDFsEMPNGT
Dz5vJwsqVBfyh+s7O6dMex5Y8reKyyI1XThd53s09x9R10MF/pVpGKh4PZM9IfD5DiTZrPSYJjiJ
u0OeO3gpOdQjOVb1+ebwJdvbcZsIU/s3+X1JiEldrc7C9bLQKZMBsN570Z/vlEiMtnk6e7wWzDcx
uVUI6w8+En4n3q98BtQrPuel9yYyj/S9ql7swrq8RxZgWt72glXG3HLQR/ZgtoiQa+hCT71ADnym
EpM9mef1K1nkKbC8FBHYbn3aSk/YrnFErKi6pD8/ulJHKrGt4RSrBnTy1T/pbnjI5rUEoW/X2AE9
U9a8i/6IxFBp/b7i0sGqKVlQ7OZUitp6bT8UOPgCzkdss8nSvGq0DXdNqJJ0wBml1rP9Dty7v3TQ
dc/V4uf7ENS7brtD5c8nSWZn7QRnq9bM+FO08Uw1fJobekt6WE2DYDFfVvXAEq2USjsj172lNSK/
m3mT3nnHya/dvgR8xujovPyy0jAX4hbBLhLOmfDiCY2TBov2FcUvkdAO3SYHuJV4yeRr6ko2bPft
kuHdOLtkShII4Pc8sNiZpgPUm4J2vHTpD3qXtWiFu8X9eoTKZwgJDqI4jG0KW7AJhzdD07kGZKA0
jOAsG9RUh9TZnpGBGNJM8LhnUFMakGpxsHZYy9c9WowGUXguilTuCBHQjMs9SP3dN8Xh04m3RoHl
IHbP3bht84jJTt3Y1bJ2SvkH+PS02D1lVp8I/B07yU41pAlxb618BtvMEdi2LLd1Xde4WtV/SKKB
s3BcvXSvbYprsGJaP538cdHnYPkxWd5u0hE199nllisVphbiVajB7PD/9vhmGT6ZkoC/j8dD8Zd2
HqOZlAFjEW/uf+MNDhrTXF8wpI6ElqadgIwePTNbmPu/EG2fgKHYv3d1u6gS27PgxKMfnvH8ia8J
XHJDSaYIGBUmhfF0C+Z2gwKJjtEy3Hydw5yRWzkHEH0NpqEHoaP4ut/idbZktuQv3p9QMVsIBo20
EaOLEl1qKlKuD+4p2UW8up5zCj1O59hzgflLNeSOoHo04Qi4HrKBA9DzoetylEb4uzoiWpyH9Nkk
DWzkKfAhD3y0vTqek5DBlbh+cXIj3+YQu66Zbb2SfHEI4bs6PnDVXSxhdbcSrIEPEltQK6fx7fHd
mu/h6IRh1SWKYNgMJsU0AQR/OmCK2PPlMDJBqdIePE2eH4uOqhMwr1kZN2PAy5AsE8zsqjMsCNJg
QcUi/I2yB7OPugRw4kpHvZkxwdTIRQ+jPmMbRF/RU3vUVdRb1e74AZ9tn2Mddq5F73CXJjG3PfOW
jwLvezAsCXn6K+EzIq+0EUnwWRZSNYDbEPoIOnGNgLQhQSL+gU1V89kJJ+30AouY0X1+Tp4hAx8F
j6VUS4+X7tOq4vcnPBimghiN1IHMTFQfXrx5IalKg5kPsohc5ouwtTSfeUApf+pTzNJXDZXunbP7
0TypOgo+cDeGeZ9GYiBeEdiYeAdTr0qoPCCnWXrAyIYOPQCY5dF7JU533NfBmTYI+/px6OW8/skj
oqDzwSBHaE25rxVSh9yIRHDDSHKVAcjI0KcF29Mw07UPj6dDZMihh8q31cgbZQE6cuweJu6dU5Bh
9CK7suV+uZTwxa/UFIxLjsC4BMmBv55H/0uUuWKcKSPI+DuoLL478rcPsbuuxt0Jyy4Tz8nt5Dbz
iHmgNsMFRuExN8tRDtWm0E/RudeKrxFc4DOQdLBGwaEhb+PtWOTd6+NsHuTDASuXg1GQUSFxSTUX
9kZGVbMiU/X1LEjxgw2p3t3sj8YlOsDmmmpfZjqo064sZBDgu6DMiLqG8wURI/BMHUsQTcz6H9P9
81r+zZOqKmndbvL4wbP0+gQTX0efisfAzTDhP3+5A9mWyG9hP/B3zDl93tNJYm41fYsuEvGNX4P1
C0naqhkS2wJJu/6YTxL72YGnB2FoR/wRNnHNG6eWYR8GcscCJBo6QGJioEWAWdGsECO3nun6OQRG
Xi1URlXl5IDLvYxU5h+Wpl3/YuGZ1wPEtQztTu4aaachwFZ6Iw5w6gDmFq5W9vQSM0YYiHZc0lf4
68rhC3FgZzJotICqBa1zoH6do4wUqY/IF9a9IVmMQTDR720bm9DTFQ+n1InHlAaZQaqlG/BDyvuU
S4cUUYCFGdh0TYSnehjBFBducFqI01THqlA5M8IbcDdT0DN0wXama1rq5ET4/BFITGWkX4nr5AJY
dbEn/V7MEyxjc06bUIo1K4ch95vVyfBgg2hogh4b7wjmsJ0Xz1tgZkj0DEugFqjMvhs8O0ZDV/Nc
IIk5Rs3hcKaHRTf8DRaOAOOmKyz7WB7tlfg6nopdPS2JLAp0qCXbANqLZwk1ACIJtmOMU/Dcnw/N
JQ0VJT7Sv47Ix5co/vNB9cYHsRIGkgV6CyfevUk/EM1uMzwv1REH2fRL5j4y2mHZlUABAHqs/mzS
gB1LEibatUvUDY5iM9HH/l0KpHHIhSLcEgRM5pHQdttiFFMnyEosrMHkCcKdkiSZbpJcKhD/xHoF
tpMWkWAPC64p5Yi4WefyTP/TRcjNLLTYiUZbMcYZViS+Iopm6zu7oJylMwCui07QsuBfImKVRW/z
qMo7w64IESR6+N+A28367oT1L7qYBemaJURY69IBQ/RP0cL0HFFL1aJlbUjeaqJOcT5KOjmeypMx
xEG7MJ3uF/djJhSjzpXy14bblzC/Ott/L5dWv3dYkgOqE5WEl3OzkTfT9nb8q6Yw3GLMLOIVa/oG
m05MCHN4D2tUvh/1a9TmT7xB9XuaikKBy61c1E84xwLLHBen4fz8E0ELuOOa4h74+KrcvnhUMt7v
foLInuH5OCnBGWhrhIb9v0oWXKEH2PZ2SSD0KKH2yYTrryAYPgtIMGwNYwAfSrlTO0zxqS3H9a7H
TP9EuLBQJG5TI5y7tNZeOCdFI7qO67x+IaDJVJvVdcwbWPH8a1c1RMUSUdtM18gYQqNy0olr7t9R
sqaDODGK+bksemAfgsl8HsjBnwKiStsLqMnwtzaiv2l4frLtTvhP+VFz5KAqfN0IgDEZkY1jyG+A
O2FHSbvMemN66aRTsfCyk9HxIdgTudIFojZzH2rtwxcpyhKFWyI+myjJh7YzZxc5XPnMp+mOd998
vPzd9uvRsNN1+YCUWyhtOJaXFnDcN98uk50vFmQWN3y6SmYlwp+fc8Hfxnh+9OqKCMLNzg4gpIVj
dt4tsLN9YeCO/MCTe/o9CcMr/YKdX90EPyzn5ToaQodmsu4ejQG5wFeliaXiEb/g+X4rySDpY6v3
1e/0LS1Eusk4xRV07xK6yoe/c7nrqm5UBtFRiLwaKzdsUKipQhEmXGss8zPtOrhmNzsziXp3r107
h9uq6KuZIc+/H2Q1mCdketkgaDyYccvwJvaF+USlPxSBy5sFJjO1o702hY9qJtFDG7cOoEy1yAvM
nSsc2L7iXUImYa8yrEjbmY3P91PjkSu9wTFhMuHQf8c5ffpCRyyjgaRoQ+FA1vCBdq12K4hcKJAh
MdFjgmmgMLD1qTNxA8woa1DPj85rVXqw6a/zLxfEggKixgctIxh9n2S9Ug0k929fsGWB9OL0URin
E0/8NymBj89pZSYcXI4DzrfnM3oMcXLZcwlC2ziTFeAXrfm2A/NMA1MPCuCQhbRlJGq/AP11KmB8
mjQzafbT0fUqWXmveobdp0AIqPXireyha3qC1EkeHMcwvHfqNav3vFfOmAbVljaf+ugYmWmCvRRz
r4UdFqpUFk5Ydbalqv/LzpYJiFrae3joAFGqBsgiiRF24SECMMXj0qyP3Un702DgZTc/82G9Vcn0
jKbZsRhusol9dqEox19sq0pnLkIH8wA9FuNJtdvwEtTx8p9oTAWjlReKt42MFdVJHrxSDyCVpxIz
ioyLgEd9+4GM+/0wpl5YbSA8eBavDm1+LuUIfL/zvvu0ydibV0Lzafn1NuaBZrkkCPxeg8M+XTWA
Oor+vttxfSUswpfBtfaWRYevXzd2mi7nTv86Ue17iMzDf7P0R7bEVho/CRJdITR7lwvLxkNPSYb+
WXMK6BzC9tszCW7xHecUhocCvKHCSw/Ub1uuvZcGq44gZzKGuc+mlEqzXndjgPZmIag4epSFBO36
j7+yWUEy3U7PJfyXCVLmygP4d0FH/gN5JiI0bGSOGARUy3gFJQI8OUxKsS86F1DNGn5Q58vflVfm
jaLXGIfvENNHhaBO1b3p10Dg+RaAdAHE/ZB6CRIap/F+8G2JFNGzpiiH0LCLp8pzmYqHoa+gA9tK
FYl7No6Vw7CqFI7pv7jK18qa30BIJrIlL+4cUXvSMJSWlhGF15f6xcIvzxDOwcW+Arhi63JJcqUp
88q1dwpSGGXUKBqR1MCi63NQhuCXUAC4nxKOOYoURIb4BfU0EEkUjXnZqgVm8Kt0Al5VasuKlxAu
UkJmN9A/JqYXEDgUg8FOMDGSl/90Le6cOyy2Xwtmc802P5+fa5p0X7uu+V9s4BTZUz2/rAGKexhZ
lSgJ0ZtXkO6qxyN15NS3Ijl42VZthOTsrIZM0tUV8au4kj+61jz0Av1tEOtirlgNZELhD496dDal
pWCpB9cmq0JHe7aDi3NszB3y1bksRRTFwzQU1um4w319Asm3iaY9y3OPdMH75B5pyi6BDc2tEZP9
nHufxM5jzWLny87n+QM4ux1nFbg+hkdza+MOToYAaq/snUbW/Qkwyd9f9bKL9PcNYGwI3EhJkO4h
eje/zIXawFldPw+j8fKqEREtNYhRctqPEScXNTJN70Flgv1X6Fy4vCevfI49r9SRQMMGe/93jLMb
RLHl/uI2jHTmE4Ggxgyi+v5fWK509Er/jwQXkFwsjV64mlC66BL5typqbXe6AZ0JyVDG/mdDUxYV
/fDGF4zlEpDGYV2dY279EvY9de45ELENaycRybzG5wptj1hmQtpgXYPChkGH5bUCMV9/OAhZslZg
M87Gl52a7qulnKdqQlxog4x8D5jb5KWOpqj0kMdY7PZ/B2OKNAmgrU+G1wiNUydE25M337MPcduV
J9d5ErezWlcw74rgAqmeK5fbi8Al5FKHNCevPz513wqZWeDjai30ZGvotSu+BL/zK5Fu1JehN1PY
57bASUat96or9tDn78dW2RDgWyBfWUxTgO0mbvKwPKXhJL9mCPLV3qClNSRi66Reeimfbs6ZTHQu
LuzGmjseKmtb2VFbQ83rcGDusBTLnTdmUkP3yGpF2MGSYaS159GJj+pD8IqZM1etbZ6gvHX9nVlS
USAs6MeDIabC4ySCYFh5qb7hj/u3Kzru6joXvzIckf86/T6LjZz7eOl+t0UJHyYUzoqnWjApTKYx
bk6a4WyLRR2/avOZzKf4VVKd9jQyb2CEtcrjwHwTxMTb3GJdlKN6ZMIcQm8ZyX0fD3ard6GVXVtQ
RFAshtD+CXXoK5x/oPGb4TIO4dhRxhN0T8QdesUC4vOduq/gbFSC3fSfCHmmE0+H5aUEzvjoJ6Cj
QGN5g8+ioxUrcguWGBv2Ol6BbUV07/qm7UkZRMvTl1PQfsMXw/YPEw0Q536jYt8B3w+yjxtKjxd4
VxPjeBiwlK1TR2K9rsKKoSRQIqKlLNkPRHAXvggQLVOGl8SKl9xov3qLfSfcJ2d2lIj4q8L/YgzG
Ns1CBNYvvS5uDC0iTkJ96aGAgbaS6NCFWE6rKE/vYVtyjS+q4+6aq0yjX5aPJX5ZE5WgZKB95zUz
lA5XNbctz0lclnFemAbKqf9ighErMYMainXPYbyRlmGYEKLoxHznuOUMJkParn5ve3HOM1uODkm6
sVej5cd+ErUNBK1ZgEz212LlI00OHtaXi1Tc5CSNT6GzRYJTSe8DKZlla54/Ef8kysMBSCfrje9z
hx6v1Dch4Gnsp/eDQeeiZzsNUGX2Yb36hkH2NTxGN+4E0DkVwWev2Jrs4tnSkULsLwPEkCtOazRj
OsGoKYOtwhk6sEKP1M7EbwXGW/BPSL+ONZNYlj7JfiwjMsH5A68cWsi+Xb8N/Vv1wucUZ6Ky5Zat
uweVmgRbt+GNeAv8+zcjSoeoeR0loBLTK8PVqvneiQ9qHZIEzNaqs1bmORBavW4sulJpHVphqGuq
ked1HIQC9iwKnNY1M8k+bXaCFtArTcT2HFj3BEYnB5obzK35zFLDtqJO2K2jQkrLpJwQOmL87Td5
zfsITN2mZA19Wvqb26mmi6gOBoN+TwS0IEk8j/NFn+JbITzlfS1xpanjfwf5rTR51xWsfKvdF6g8
giA74KlB15JpicFvTrXK2FuuZk/9r9XYuLlN73PerBfl99GBxxkpE5zA2yt9idkAwLyLX74jzQZv
BL3rgzvqEypUCSvl5KvQdy+1JKwOxP7D0JXIllCUwCqKlHq1chvinSWxpy/GSH++sJScWmaKLppD
/Wz5Vnklie+aZsceaIxmKQQCuuzi2Te4nFCpiEDa39DfZIu1foObGsoWkO1S3KyzJCDzWsel1f0q
aMw5YK/+45OVd6xY5CU42YpFbP+iu9dWdwz5wik1HPfXS5xcDMYKp1FHTByIeEz7CLVdwQc/gO8E
1L6Vgz2o1jBQ6eLWfz6aa00GVTKFAAzIqn1Pwb4+L2l0I+P3xfoYQeXgCBM491GTvNm97ndt40TF
pF99cLdoOf2nuSxUOZEhN+YvF4L9Z0qDyMVpRAI3jilkNF5xB7V8gEc3a8+WPS4+iVV39XlvNBen
0+yi5/Mw+39a1iiCyTZGfjXypPYvrMOG9CXYTpOLqH7x/dZf3igT0azI+2tk1Q6YRJ2sAhrrqQIA
gOn49Wsm1EqFZ1siABF1C+bhGpnwj9lRT7OUicq65x2r217VwCLlE1opEueqdzqZMUtTW5NYjpNB
gZQQxjkVIQR2+lae4DwnieXP1CHUQN4ORqPKkfxBmkyp5/5kVkyI1Rep8SWJZqShO57Gatmj0ime
yTB+KIhJn2g0tYt2ijRKg/DtNBOiEHHGLIPOtdpafjVRKlkB2y2ba+MMbKxDsAt7vehSx/7JWfIZ
FdRxucULiKwUlbw8Lxf7dWK26DVUGX1aYQr+lvyiM+uhaNRuSmaJqWBWFUKD7YrwAbEhTWOHFq5g
SbtlZtV795uen7v0RRWdob9AsYNJhuP9FjnsrhMizAPa18Pgfp+2p0TKniaE/qSGGtucpyZBoaEc
LmTJ3O0YXo7gWAVU9nr5QmSnJPhpdum6KmiHxuFIxg4ZWvA9XEH8TZvf6asqgzD4rYkMxYADbKxI
CsPvoFv7pvtO0zkK28s43ThN+wa1OSTbcext5riUhkhKrSssao443ORhLJxMIyrpFCkd5e692MUO
kdFB0mNWqzjkim67PX3Lpz/8scb1PdSHVHruNLqJm3+bImDUSaIaH8dxHj3gOgGbF4YuEsCEZi1V
yff5o6HggX74WOrfIG/MyoAF6W4ReOH0ddQvK35ttxLyOiMKXiGLmh5Q0+TzEyLPXmDrh1J1A9ys
XTEEiC3G9uuP2X0tryzXn0yrW2ZTcTHi3H66Pu9Hz5bfKOE+khfh90whTKpAABVJJRtGLmV4nZfg
QW3NCx/G/DWAjZ+ExReomXInjpHOlelA2wXrKFnNeZXINxDe+QAtjYhcPeIMkROfaTMl7c1kd3OH
zUKRimbuoUaafdycn1e64Zn5QBVGOC7QnnGT4NmSHEH8y7Ljcw5DBQlyTeqSmvy7bIbsJyhl5GYR
OH8176ezt6zMmd2WYS8riYoEwOczzhKL7WW8uKMpbVN/Dd0CJmEI87/BaxUKE0BbVFlSLyvzdXJx
uJtk/K8VA85XHwe+igrYrbwkBszenM376yLjyDeEfokfwmjBuxek9GNNoTmgfhrXKbEelg8e4zbD
Rd1Ee2sq5cwmuLuHMnoOW+KHSJIpXSG7AcktsZ0gEA3wp6N/3uE242e4hrh7OlnMDMKnbKI32E1J
hLskOnO66HaMiT8UXoD9pnF+coU8Q29dpGYxb0xhCktL/V/Ae9m/08exGFk39H3B3yZLBGZ/Kud4
ETJ53P8B4+a1NQkfRtz30m8F7x/uBbhnogIum1BwWumztiwzgW94yDb7EgfdsdIzjEXsV09TPngO
bVud+Gp/7Bt26zWMjzR0sIYRXYufApiyUpz7lEev5lAXNzULm14odmmZJV7oTXBtbl9Fxim7K3Bb
kX2Mp189yBqy2M2YPBt1XxlW5ZRq58jIkGgJZt7qQMxOqjWHwZujDFJPCB1auQvRKHGSna6hPkQZ
5PZBI0jZQdGdwGN6AglB3YTp0OgT4WEIDkO2JG3b4Q6Nl7BrIob3nH0o+BAQ7KhYCzoKEH0fRE1A
ns3cW+wIYmHlzHTL/QM3+iPVaX0DkHx6EAqt0MqBnE86/MZXzFjwCFQoS0XsjTYkDVlWpqRo39nh
/IWjgJq+rxesB4z51LKk2idJ1f14t8E8CpUrM0c3uhrpDUjaMCZj9mqDZPw1tQoIDfRr5zOlpDAb
Cwqt9eyEuOqAWVyel4cRRqQsQ7H99RoLvMVcWHn1xdTvo+5Daz++BrtEMAz2Q5G43yLO043KGufK
D4r+F6Sso1UJtjV8UlUl9vRaYFJxe3V0V8nrm4HlBbZRn+nDj5XbUVWXgF1CIyO1rpUOaCnnSI0m
Crm293PzpN2XHzliy71PoH8y97GuJmOa4q986Bi6lEYhggcmBeiceSBUwnAq1VKJcLemkv03kSbn
/GxesnrA+cvwO0JMAsAuVMpmVhWYIDZzsEEyqSKQuUureeNOiNqwRJNP+6PMDOAsJYFZGVbIutXJ
LNOdn49jDokywdCghL0HVTSDyiSyya8I4nXb2cG082K31DjmL87/Y8ftD+ofkFF9cw1ehrY6GjfS
u5P98x4P0+NtK1Ms/oKu4je2RebCJmJhw+0KmHdsgqAv6yqKk4UEZr+RqUT3NnyGkR2JcTmRxhC8
iVRbOlUIHQ2oaXPwM9ga044lLd5Y/9lLjmwWVuqJg/VPLb1aybUGUz/p18GUheq1n+Q9lx/jgH5o
gNXPcBeRVH1jCLzJJLJHf8hx8xIEqGzZlJSjF3A9i/n1t/UIE1MRZC1UNMuffwiAymyl+rdGH78z
5EmDW2YAQxrdwXWbgj3DVqS46Zme3QIlVZ3fChbr68LY+ZpfLnYMbybf+9BepXMN2ifVdYWgZI7d
ZXUd15sF2PrZN0gFX00ILZJfBJltjKJN84dWO0JtLHMio3OE10QYwliNBJiYsccIc1qFm/Mh++YR
rz1IetbaWKZFBB05WSHTdSW1Kq4h7/XWQZwKrpgAGJhdjeaIjl5L446jTc4+pCacOf5inwjeFSMj
bIRhXkNZRogab7txk3wav1yPvVB7e7SdquiO0exmgEFuo64QdR0ob/lcXaaX3HTRRchySmtpHJep
kqAZHqKcPjWV5lVzOGgP/NTG1QV8HMfZu41C36OAZUcmcOD0ONwvXxp3tCvYRnAf9DIhTaatHgvy
H2nh452BmMxelggb5Em3zhnisDKsS0ZaiEfcucfHzlnBL8Y/TXglLkPJnFOqaX5L7sBMBUBmg0V0
gnbVFk7a+h/xtKaQMOWAzTnq8ucpVXLYXyuH47EwQfc1NWJ0SQI6GHWIJ56iT845gQChTNHrlDGe
3SnYI1+13Wrc443dAVxvHUKvJmCzKCMQyJxV958RX6t1JSUXtsr5O1gZRVzXeWSzNeaEh6ftMmWl
5bDFwXwyWvL+42fwB8jQCd7W2rvec+IOmuFIVboqsY2r/+EeLGtCVwPPjjMrN8R9H09SuHYOT+lS
OzrJr7dK4NyRrwE0El5lfkWRMvzphNs6m8++7vvsx64x2NeASL001h0hbaHul0YC+6hPl5bvvrCE
iI5qvNSBA6RhaPk6vRQKaFwzCjnBR1jsRlupCaBQNeK8YJlMUcoEkp9uBkafpoErw/mS/fgnE+hr
148OABgsSl3MhJkBMggfWAs/JhzBD7a5vrwHqqt5hRAIKU9qgygEN+h+VvwWILzig64QX0Wbo4Ol
IJLnmIMaUO7ivRprx4GZiuyhgYKqt+Ta0rYwH/0/a6HzDv2P48jzAbW1ChLTsx8m2kTCW2bQFiBg
JvIXzhxioW+hfx3Yo3jL8L2gCzlV03EB1FP8p50EwA58fNkziNQX3KEclvY+D/rR2zSrrY/Nc0j7
7xzotLcI3ONTM8AlNu9DQIAqSLUD0S9M32ltH6IuHpX2IreMYW5oSx+khA6JYc1UhWC04fV5uYQQ
g+yxavdGnN73zhDoxu3NfQT7fnMWtZQPeVsEPStBclOpAhXQjlWsDkwKUUrTn44eCLiQkXPuy4A3
mtTJf2+0IZYZdphfg/fDUWFNhBfwillR7bunPk2iPI6F8/ki/lEEtsS1UMzkKiDw2EB/EzdceTne
F0ORnP7K2gVCd/FTPBLhmTgiiLt7HdOLEZPu71LqAjt6kLVwfcSxiLvODHchcM+nuxC9gLeYUVfm
QlmNGcNy3MBmq7NnNhUpccdQaZAJSSyuee3LanS8+WrS/orS3bz0iuZHt7JrPZ/VLIJEw+w6+1iS
vvq+og6JXyuOv52FxxXMUiKwjXnH/b9BMTei0h32zrGpmbN+G+5QVtaMjaP6XUhNiIGBWEJZd/bt
87Hth0XIbKjNHgGioWb0NK/ug5/YpYgHQyfsubsORoEeqJCVtC4nhPUJj279PrUVYiJ4Uhmhhhof
pQPIXqRNSwNkmsZlL+APvKQ34oft7Q7U8pDLN1lf2QrSkRPBepw29iAlAXMjRXiDGbm1/vWHJEmJ
WcgsnyWVv17JR7tKFFioiCecRUqi5UycEIHZAraAKzn0wdjOQegWgJ8OdD/dZq1Ak/LHU1xqAKsE
+JeJzWBZ6icf0htuRGnEl0NlCeMnpemfU2LU6qyUSdAMyurnj0/ef7WEiHTHuvPXBa9cqfkKuEbY
pDjVN1TfcbQJlnLRh2DLiJ6ZGkLV2IeRo+IjG/wEbz/plknrFaiffEiCwBmJ11i+MfKJTRhhkU4E
qPRKSpRVQAyB3dQzRoUtfLUbbcI8t6zOPi70z+PwaZ4GiuqP6KFHAuEsMgVTqTNj+cwMr/IKCjbD
zRjAcSYOjvhb/co5qZujD4yYyyLcJJJJ8Ea9JX9NBCgNjNFeMnAe6FwcCdHorwXHkQYHXUtgPyex
p4Rh7QwnTdfj6/CZaLBQHC/3lh4qdh1QJ9gXs5NuaC+q2DQShBiNrFljzJjuJ3HjLaxB7egXabTs
X5W4b1rzRM1cE/4c6LG501sXaLMcYLepI2lsG9DBZS95zB2VmuaBSgQZKHVIc4ZtkE6VdSSNMl6d
Lulg/Dk4AwrE6phZudXuAE2m9FOtKbqBi4yVlnqzuTH7Y3C3C4IKugNJi4197vPqduAcdp1t4rh4
zwr2j4L/PdhXkv7sa4c0bnCZWTJ0ydC0LK8w6LNVwHE+ix0yuyvEWxzOrO5Ns9eE6/pJszxyuyfO
5Bh+szxZeuNQ1go0V5eBpaGQPfSpxgBUXG9EEGA8p3SqrLG7+S3qPGuIvBunDuMWYoJLMj/LrPAJ
d4UhRs/170OGoBfD2L/T7si6/uNzKSXybR7q+QJYIrzIeno8i00YR6c6b+Ce14TK1JlRnS2IxA4/
mWpM3I0xbZ24I4L3dv1gYd4vrxPHBlsgloSP/RDbgiyx12cbz+t0sNgkOl5b/cVkRUEasY0d4Q24
Cg/WIXNk7GB+9EZ0YuI4Fmg4G2ZfrYyO8CgTfhqihP/Vu2if/v1Y/MVoreFgFArBbXAz4zBM3n13
qXV0CjxBjZNIb6RiuNRAsLiW/B7QYjl9ZKNF/n74hLYz6LFSRpfySHTHixeL5NdE5/vYcRSSW6jK
HVdHD6nBlGjdDnrRZAcw8FhEmO25TtPodxhZxXcsqHFEMrbW2Jq44mRxqVzVfRDvd2VGhknKa5Di
y+b22Nb71p0pPferQdcnIRW5oO4jItELtSwHuDSwfbyhKv3iHqoJ67uT5QZSGe3BvUYGrsgchuQ7
wXZSQRZQEAVg7f30EDpRPeOd4pdEZkxnJVMg3xasrDXWWS+iP/quv55PH1qq0t13WR4iuKd3OP44
etsRnXKrnzxk9h55+GJ1OxaGL3FMNGowgDMmb5e4SdNvLH/VdAkXrMOa59/d7uZUMlKbhWz/dpiU
MA45cvj+JEgSML3wHjrO8e6WJWKE1r5YL2ae0rTUacZG2rr8wlZk1mQzFZ2z+PLY+eL5p0dQvQL3
LXV/9zSwRUcLWydKiKadMssFlRnAOMaUSrF+ZCtXa6EfDIe6UcDSMo6W2JuKyayhfhjvjd3tTcbY
vi7CIpIifZ+fai5I24XqceFunP0sVHHlyhumCqX8QE6w7m9B70BLWYQ5w0pOhkyo4u02KtaDduyH
Jr4ECE4tuyIhBgS6B3YmnzYA+Gpms7MmOWa18eWtc3C99EpxlJ6d8+9/y2dpngyjjYM/dahmYtli
4XMWpMVGxIpW3A6ktidixUb9aqBEO7q41vk4f+i+EUyf52r/VxVsGHri4tD8US80Lrf44Tu9CScI
VTCo0OBLa9prY+cSkeFV2b/Ecz/k9wb5iYY0myAlsHMYh2CLIh3DDjtRqOPc+8LOGuyA+UO+qXj5
JZK/kKIL3lmMXNU8BoBRKELWpriNe7LXq9q04IIzOk0ZnOirYCC7pX14R2spT25Y0YNfuRHChQOl
PEc+TaaSFPoNl0oYTZH3E3p/dLuO4DargE5Csw7eCPr0YIYfxZUPAagQGsiNyzklxPvlDvaaBf0j
2Trnpiv/KN8KOnTomwFe6W2SFKkU9fMoWN8RWMfObDUrL7XMMNki0FTAlrRF+liXK0WtdEcAd6rg
0S17KGH3KgtUsFiS0/xmzv4Bb4QHyoa6Q5EORhPjKCVHBoxmufxFXT9nRqY2ybMhmAndwHdpiW8/
m8SVc8CMAbkJVdQXMfk3von1D/U2IX2GlMerakr32RGStvpWmGLZNNlMuzTKzttN0KWg6Dvd6S5r
q+QOe/F7ZGTkdJFHFgwiwFIf9rxip6DX3xreYXpt5gBRkHLgXa0wDEmvAlNxV8kne76BGtQ27WoU
lh/a+5CwrrfV3DjXUda2V7t32kwBNwvZo/mcbORL3wuyP7JsrYj+ZyoIrTzpg2ajwASagyDFA6MJ
E1F0fxEjjdLu51+E+SzKHoa0MTLMzIYGacSybhcnJKms1JraK0trPtPESmHt7xjy64ys+yr+2aWa
VWZ6p88tnaRpFgkhYF9fln09DfQiKeAlLTY1u1aWwRE1h2TrQ4Q5bspwaWV4hR+sG6Tj2aV3OShk
W/KZt4rrt9omCYGqj1Oi19FEVblOITjJBwa3L1mrmIxHWlDVjRHbkmAOzM0xCzLOvBAO9zzJ3my2
WReE3kwTFfbRBdhVc1NEIVQ5gRabgD0rerLjTR8B+GJwZ88vXWLmd/8i6we3tvGm6o6ateM6sjbp
Jftj7vRTnYrabZdmkhhNEe6qUWbqfHYBTB/rZJQsBBDxIgDWukF5rLpiz2Kf+fVHyDryhPJqlTho
MqSVhm66JVH0WwCfmUs/fkkD1BnMrwuH7pasxiIcRnii1h5gbLP2oIwkwDcBEklnXjY3Q9fUV2Wb
y5AMOEoVcN8K5AIi5sIAkpX6BbO7XGiCJrSGsXIUKQ5kPc7L/F1Pw+qKP7m2ddLEsa2NXfOKkBFc
f/UxF67Hckv+APgxT2C/JYd+7DPxO9NO5FRerkPKVDGYqxobB0Cy3AT7lW8i6SKS+dhi30A5WYeN
n21C7SXW7cvcndxUhGjAdtTq4ZImRjD4gOO/azHPTj+nH9yc39fLyKDUjGLM3zaZ5JaRriGWOGTr
putgs1EWu+dwnG1nr0T1eQ4t1l02pC9pMhp686Mi6vJtmqHscfrSYAVIeAXOLCnmjdJJUVQyhFZq
5thify7Bz4F6YP5LiAAYKSrFzZGjY5yoHn/ZvRsgDvNAF/XX6udxV6I5qHATafGFLyqgH3OtyB83
1i/g5Cf3e+zTXwOVWHfvFyGOXoqMBCz7QYqX1Lah6j60paRWkquwmuS+qByeEc4cD4rWZzHPY2T0
ruY4OYJh4sHVJlUXnlMa2PyNqMnpD941EqieSmUsK0UU2pLuZUQOtLkqM5701dQodBk+pwGPxFvW
DE1dUaEZKVIU4C4gZ39bdu9JJI/ZC9BboGtodpHw4kwN9wsLcGFNpbf+geByykFgkOdjP3HKWX2J
LmXh/VeSR7Rvm5T0r7ChBOkk1EXzY2qTWqmTA9ccw6PXIk86vlEPsfsfeig2wRe6aNZTqWPqxMXY
FqDCN1IN7KLRfFRx216iu9F3NZEAc7XR6YO7HUPkaKmsSDUh33dawAsBEc8SGj8UiNHEA/D5eRwK
4RJ6sbNKebN5sPqPioB/QTrswXR+h/7L8uzAgxcDO+izcjR8U+pjLQHxC8fwFEibHTZxkpovaAqp
4cKXqPblBFR1b7EBaSzbSnGuX1Mo48YplXoOXl33K7DhbRGVLxEwkHN35MNFKsMlWcEA1Jt3agPe
9uWOx9bA7ApAWOxF8Bo1YI1mrF8uOagMlsKoBD+vle4oCCJ0R/xcPPGGIYG6VN7L6Gbuukgj0xDF
gFsHK+1owS5IR43d6YuAy2riwY2jF2gVc1GJfQ71sDaKqr8dq/d9humJ3a7YdZiL6/+rtL3e9XqE
wFsP3kjjBg3dkoAMQkUPhU52/y85tAQ3YmDzbX0yY+tVnFiHRJ48Ge/3ERKqEJPWIqQzdCYMjKMI
+/m4jv2bGwg1uPIRYc5H3ek3Wy42CDz+FEmC+n6Uhhcux/Lbv40fJHUomqbGSou9+il12reAyVVD
aoVigZ7ShUd5To0An0JQG89JtoV1lXwCRX639ItRqG6DRA34PuUXOEn3xCmayFJPaKK/B8F8xqzQ
ZjKL2WxK5cDC5tIYMOYb4GWEfk7XMeegbJ8ui5ti0Gops6nly5tOI74djkuxB6kUA0vY21wgt7IO
uSXHpOYlBPAQa3dCaRBtWCH5Zz6idgXkVCc3Fu/rO0+Xb/KjRNIqAQciN0qhccsMsYaeH0gSl0FS
50MKMncWX87VR9dL8Pqd7NV3PifSRFksJrDdZ0FiUpAJkXHi6/aC/UeSutAT8khesNgWI1Hm6ri8
0KaYGq1gCc/XAahOhSKRfnT5GNswYiEAIbN76sxCsV0KqG+YQgvZCQmOrN7TGrDQikof9/dbF4YS
nXX7LXv0pGEP3WHKkhqUvbqP/a+ZZvCgJT5iZUZrc3YUVMKyezsrvt0nuWIZOo2fCk/w4ZK+/mkl
eMGxP/tKsLpCpB4tTvVy0JP0rAr0+cuktX4lfWz3XGJYNhNTII4cYgmVkAEss7Ae8EmLDaEwSl3c
8fyCFfybCM+X8Mz6T+QPCgVYPGq6CmI3FHkTA/jzYdFgDEWvGXdLrXmbeoMVpCVNetXXtb5Rkban
zHghRMdzqEwaukH0DiOWovxVe1wi6gtxRRISqEzo7jTa0tUcf2LMXIk2W5CiwDXzWk4blg+nkglo
H9A6n/fuPua3Zab4SJ2S6/SUf0MrNc7L6RhUS6WESsbMY5PlDWmslzwmM0by0ENx/BD52yVqfKvG
uBqZXTWpnTUWOsupnYJ5K0nD9wfvYXyIXrggkvv7EJu7qk3ltMlWth6HPpCV6e8YvlUcYkvKIi/y
tlRxDkcHjInENSiXo8E5DiVzusU6tbmU4GIa3xMFa/BpuEQEXSEpAwlC0hNllzcEtgDb70jCf5pa
JiIr/Gv1vOaQqHZNfqsjB2WBc+OCaoZgd9x8Ufw9j+gp2/twqfOa+yifa2Etw21jcoytFQBZ/koT
aQpeiNcSIQGXFT5N2p5EtSntJrf9gowknDKPrdT/nn44QvUgnyn47QcA/+8XQijOaq6nNr29crwr
oxWdzHEdkfSipGlwcdPTjCUK7Mxt485/YM6Q5f+DOXDani7/KQlTUl3O0vVrhpWiXR8W74mHQWIZ
ZxCjEThbIhv1p66yEJOE4vUEDG5IK5arjdlzWuGAzFHpauqmG2PoNFJID/Xvi5hiokIL7KAPlvZu
FEB1wkxEY/zjJYcj+DH2fsneCp+sSmeqCXAmwl/5qrRorJqzu1TwDBRPK1JXQl+Dv/s7IufyR1BL
ZdqW35aDxRuSJQ9mq1I9vOoJ8w4hr59wipYy7zksh/bTgyXYLw2a13D4uw5qBMpMHujh1/1fvtNB
wIi2ogGvPMuUWXNkGYncP+QPmBeOMYnEJ4+J4jrALqEYBRhzFQG49GcqfZz+E79F/ynNhRI9FZKl
dQxtwe9B36DTLNi6RA6HVj3tMJ7mYOCJqWDYSEcDIxpynk3B7kQ1OGQoPJf5kOb8fI6uNhyM36kp
wZvWJp9TXMPtEHeuH3GxOO6yMxzXWAh71C4n0iqc9zZ+7+UzXUIkf46JiZd10waZ/sl6Znj0egAf
gAx/cHaeBAeMxSPQdY0tIYGfAvj3M8R4ONrXQ8znnLxPUlqq6Fl1YWTDqnoY0B+HEnGLsTFhXZZB
Watcsk7A04hmT0aXQWMVbcPBieeaLrLhOnowCYjtA0bBojXmI2xEw+6OZ6VSnqSwxu1hoj1nt1+A
DKly/i7v84r79i5ud8JGFN5obM0WwUBdaMqwdAgNHdm65hRaoSTIQy/VPyQI+kmPpK9mZMTn8ymc
2N1YtTd0vqMcqWHubFUvL7s3Fsqog3hlF19ZYAGXTNBTM8+PQWAA9sg7xH7AkbonZMR/PDR1U0xz
ARBqV6HPPxPB3GaAof1qP87h2tN7U9AFTxTZ1Z4z5ilo5UdNu8H8DjxPre1mSMWrA8FFSKbpEGPW
L5XQJ9T3CErxNX+HcitskEXQQI4VodKhh24gDFu6w/bbbmrUcPzmxgoOqP+dkBmAQfKxHuYzUJ77
6g29ijVEvH+kuNKIQ8PI+HIa5heUztCHOY35T86WzkBG/uNluGHdko9cLieKRtc8MT9wlQx3wapY
dKOs/UTbRzNxAaACC70NF9zaYg045sYh+df9MtW3EC2qHDIj+m2DrS2LtkAwp+vwAcAULpGS4cFr
ByqmTwadWcfWsHSvtCA5WznlGXApwAjOWUp6TQfJa5ag+w9xs7qKSNJokWxLvkDQzko6GGizSUP5
idFKcKdUCmDZXrkNp17Hhm4rZL0oef0gUPqo1JREmS6/TQIvM4TKwkVLs3JmVg9TiTTmJ9/d9y1O
DoklQckiIVSJk6NF6SfTHMBlZp1K3pT62FW75ROpkn8lY97JA4J8cRO7VBzvuTW1F6CGsk5pzNsn
EsMvEZS3NnBFZYrehxropqQAxtYUxgdpBS0fBv7Hc/c9pJAcgi2m2DY8tAKa553mC8NlNRUgpfdR
vjSAUKAkSEdMiv6rafdk2fgXUe9Q6yZiiA3a+0UsebmmxHJOj+osUZwlMx68ys3x2vjK1GH8grsp
cmreUiE3xNJzaTK55858AoqaCH297/RelDNowd/crJ9L06fNIlsds5ZEDc7QTXHcoeKW2aP/naGl
92xV1qN67Ga8psbMh4rcEBxtl7GIctXZxeeCmVUuyeKJVbRs9FbWwPl0enVAC7OIZANpMV+1xTtC
YQRqME8y73TUrBCcpb8X/p4VD7rIoxt4rrFi01G3+hd+S+ImlvRiS9ZnfOU0EEpZTNjvWn6ZSUSj
AyO3lvJ1XtwcYC/hAqtnjwfg6FYns6sAtkpU7E9nFfCGXd+EI5EO2hD7pyELlRFDmjI/V+BKcdyY
ZgTX9xcoLTHzALui06DZ2hl0r8Cef3L1YFzmWA33ZH38XC0xukkJ5uCFa5iLnjIABWi2hO0Q8Vk3
c1e1qT9X4pXyQC8WN0Xusm3VxveQIersUmj7LGfoFpgH9hs/CYXzpZNoR4Dp0SRs+7E31RH+H0XY
6tsWoF8k0rRc6Ca6ZVi+48Ito1TtSwLT3TxrgjSHktDAPb3A544qT6/VMyNOY5mBfL8llaTGo9WY
cJkBnEVg7qHfM5gcKTueK8ubbHVipKI9nEbZE2qR2gFkWksvgjDBNR+IgH0zS3B99vIC/lNxuEZ3
yfEpZ43eISHq7vkZMp/WspAieKW1IdwSWnObUJl4tUeBCuFA9bRPObPj7jN9D449X9TI4sVTJuY3
0lWLvJSGgyNxn4hz1QcDpGntJPS0DM+AqHcJs967UkkLbdcydCtnpLz+Hnmh0gvv8seW7ClZqee7
htCPGNglHVYNsYoiw3Ak7MH2PO+QV7ISSKvPIgqiip3+OCoEwhQlE5TMbsIRXnHRX9u/vJfBNb8C
leZPpxqapDaaRu4yYx5cDVrIg2MC+eUaBkM+N1BfkHxv+DnA++SKQFmNltknKhA7xL6/RcQ1i5Ss
Y1lComN7puCWZ24mmTwt8PtNB95mC+D1w8YKaBfYv6a5JvrYSzbiY3C7QixH/P9rntfFq9W15iMb
nYsIdhsdGN/2zaimNpHLDDPtTA+KVHYPpygWp1rdwTEWEkpCzEVNlnGi4w3G6J97044AbBXwbQuG
mOW9wyFds+CVhKt4HvNkz/akZ6UhmljeU9y85kjkbvBaA71YUyNvZGNnWaB2slD98giOeyHGTA26
hBXd54KUimcCEvKKMxiS++kaC8Ah2JLOSOHw9oXDC6ONl/HoMsxiMZk7SU/UKOVNDjf8jeJM9IDu
IjDe6IX6dqwJB1IKaKH7CrpTvMPBTGnQPwZd0p0yahPGK9fnorq5nWlCb8nvCWaTY1YXJNvfyrpx
nuP6rvLo/iSOXW/h76D7hYJtxk5tu1mRs7xDgDCK6smIYTyDGKqPaA7GEE+VSl4ru+3JcDJzcXLp
vWy+s78NBpFFUGeiQoCNMJpIJoCpeGLsHoVoROt8f6plRv/KNgO0bqvs/gwcOo7lTtU4JpehkR/6
puvr1qXqPDPXx4HjMAiKNDIm04xcL75IuKJfJTCx0l4ERECAcbWG9RU91/1IZyKdVAHSJjgXRU/6
hBGwyZvcAIwUAZxq9l7mHwHIlcCB+Y9CgrVHPqy7Wk9BfMipgu8rJYnoB592wmQCIiv7fd8ojDqf
MoUFoM0iyH74nl3iSDt0a6/NVjWgPmVXuoeTfkpvZumX5AfHKYd9Un7uGma+s7B4wSIIAXNcHy/7
7VTb9DDmXH12hyR/Q22u0633+lhuaGruqeBm3vj380sGfD5yuBmsYoztv4IapuWM6CcRiI9OfCQi
XGKlruKhauGCbgOPlYoIzjFcuKHx4DRaDVC/cPyo07ZOeJ0r4CW68j+TTSbEidkf1aDWLdP6MWwl
tq6ddjtVgG1jUSuVBbEpiWcFyw/HtrbAWhQSjGZ/wzq1jAkLi4XhQfCcdrCeRQsz7W8inq88WPpw
HY/B30zQSLn1papyhRToTfQ2W213X66KCBgjsDI3SU0b6GaTWYMlUMIjFjNr4C8jN1ckslPpyqw1
1oP15LMf+BDtABlJto0FUOgwHKTqjtrRs8Phviwk2dWheTGlZOOSbKXiB/XgtOgNdViWiAPOEH3G
fZlo7iQOLLHOLXz03fv1UPWRN2fLQkoZio8xhSHBCNve+8VcIN5X4KQQ8WMmtApp1yyuLoK1W1//
djowl+l1QiUU2xIXAO/M2xLLx4MLiAsaDfQCsI02gz/BRgr9JoL+hfpib4Y9qzkrmAahPwtQwCj8
37V2arpu1OtXS06GlV4Qx4NfBwsR2WYdnfuhQnzeIRqllobYQhPu9OUS6EtxcGuWP1eHyGaKwP3u
umUifqNxO4d2ezTa7yHWsaki6UtCLNzbszy5QJdTWOhW8upw/Km8aNI427O/aElWElFpnkfpMtoT
bSpxEw0xYbxZiBlI6eM9e+YrMOuWVMWZS9SBpnhSFHzW9T3bc0kF3aUurnOX/GR1dZGfOhG4bYbm
uLVOxZqKRNeRASPYzmWJFphO47q8TtGcT4u9D6+thijZ4uXwRdqK8n58K3cDDM1FMgnLALv2o6Ed
CWhUgpBktMf86ilKz9cCgcnEZV0yOaGe8ygrDf2axZv+D/0pv9cRVpTqjib/NCk2uMrhXGRmK6Pl
QTpUZWJj3K052FxHj28sF20HXJYJRTuFy0bQ8PPfTtZOqUxmxf8KGFoZHCBUoAYaClAq8DvU0PXI
l1+b44Lt7q0SR97aO8cjcxUt4/XvH0daiFnhE/g3+tPznRk5+RJIQLABpwS+YPADjgQiSbVWqTys
uR2rEqsdozsYxzRBR5gZgAe1IJCl2KxCxX/KD+BbC178cKzDe4gbxE4wziAxRuho0StJUTN/1Fqu
PP05mbS7ZJdM7hIVja+KNBtBR9ezRScYlpQRfzDW/gK/T0dpHzMOjB2+P7PmWSq8+F8ZIs1XIZbC
5/qJijvwYt5S4SvXAsQHOGKK0ePYLgxNoNOch0JIlvNxli9FXJE00O/Ja6RYi2gAi1mEn/ZlRXZH
9Vglv0s30n5zbL9D4xNnlRIqRsd84r4ufx+HROEJxIFmi5orKR7Hyx5RXkZ8Hl3vOX66FFrqn+CU
MzZ5OjmmDagZmKdfZppHfIS/otcMkbHpqk4DVHtH7WPI1oi63FqQRe9ZZU4owJR9aTcvCMcB9ZTm
Wc7crsRdCapchvVdYSrsBW9UgDcfgAlv+Wr4TnErCjq/iWTsqe5uE8Xe8MRs0VQvrkATS+XMu1fA
CQ7ctzzHFAjj7eqoX0vDSLhPfs2ua7pU8S+X2WqnDz1WRJM8xkJtDfZMFqaUkHkEOepsfiGLT18i
9GBVkzKejWMp6bzk8c9nG7Iw1hitBUMwsrBbSqEG1YHz25UaHfTb7YI/N20zTdG9DX6tujCxiYKx
JlLSJ1JxFjoniWs/pzIGCPtDQHl/po1neAjMFpBDHWFW26+Ubk9R5JmB2iO1warmJlQDf0HRL6CQ
yiD0jURBuFHgPCW2nwiqWVLdWvlB5x1I+qSjVeWAloeyLsSm5q3nMWslL1i1PzDaKoyrrW8Uvbn5
r73xUw47x93rB3ZUP/l+9ChgwqHQnSaHHSNZVTulXW2Z04F/QtpynZBuW1/z4WcpraVxhsR4i9p+
Jl305YUTqF7nctUi4oztf9LLAX1Roubfal1ckZD8tqR+L1J5RjbxFt59dRlnjpssTYKDcNNNJ+Db
AlECbk9VGSbpPPedUmXoQ5hN3aVqSaIBopMQQ1k14IdS1F4RdY/ZWanwsBKYR/1grklzUWXOK8wO
KcPXirGIXR49VGnpg45tCwQZ3Rfqept1AaIVlWuVBJv/4L2WcuQC4Vpe78VPF6/aHnFysbSK7kJA
JO60VHJ0olVNCdgSwSGy61Eqqzmy72kVbIBfr3xWRPXNsjkycXESrZfc/sZP7eL58ZajJ0DSty4S
MViC2XOglaK86WnXCHalvkBSYFcUVzUwPYsOPxmz9phWCdf2LwefVR/V56VJB0sfkkgEfWg0C8Ox
znPhxPA9o1YehE7W2OyUYsPV5MYFWn0Dt0FMkaEUkYKwPWuT5J5F0d8HYhncVihtMohsYxFn1yIb
dtoPo5yNGvxSIpX6lWfhaccpZEZYrBHYEnst8xSAhkTUY8Zt3/a57IxGjTpBsqSwa0/prVLzckbv
phJMAbKggTzYcS1gtcBH3+BwJox9FXsKaDdO+MUmiAt7TW6Kmcn6vaVL0yv0wanLevG3N0z6+067
wcDXVO2rAqc/Dd8TzF0fksDf071lMEZKItZpRCGF4YtpjWDwrcnxs81Uq8C/umSSWQsNMSjmpv/8
ErkethOOi8kIffdB7+27rgPWd8nkVU+Q6Q1HJzGgDDvKBgF2TYXjZdpc9/gk2RuyGBAzZhaLPxOQ
GDnajIkbRW1a57uhOMctlMo0Br3ZroE+HziV56TpOnFA82lg6ng8MJv6Ulx2GweTreVc4ld1DHv8
r7c1wrdexmS1zd0/BnOU0oxNVJBZ/eEMrQh+rSI+oOMA49s7prvw+1DeDmJKaobbbbPhDYIE/alI
vqQFeicSZzsDiiWulI+hLWmvibbwGhmFBiaU9Esqu56GsysWh3CqmdHND33G4aBvueFrY7WJnUY6
/3i+moatsK+86N8rpy5EeTNHRJsRf7qclLaCl4Mev1LxdSGcO+HDdj3v2LX/My5DOKuqYbOCwZrC
YV7mpyndhHisfPeq5EyEx7ueZdf3r8KTSxFfX2UY3oEicrUafIT5qkAll0XE1alAlEvL0pkdjU4d
mCbuLl8o9QlfhDXyk7BglQ3DQXqduZSumrY75lN9Ei62gbauQIpfw9Vc5b7QtBizRqt2gqAk+vbb
dlSxOpL+uJGMt/y6UxA4vjChaSG/HhEiwZUu+9gxzZ+hm94FOH9cSzsd21dAQMi7UNklVhlx+tes
IRTlaeX0LcpOZcrDXAt6iHV556fQBBpISV/tSVujQMQd/IvgWzMVTbzrSRuMFkDhHDayI1G3l0zV
p6FCBIP8k19GTMGlarfGJrE/ftmHplCCHL5w3rmrss0c9189NKoh+Vv8mTYFxw67bS2nt2/v3aVo
z1GFypIpPOCGpUq0QD70oseAcYFTNqaC2chexZY1eV3XuHkdFK8Ca7ImWdnJX36DeghjLZSxEcyH
O1KutymnEHNovAU2GR4BIHMT4hODT2p8s3dTDZvYZAL5ixHnYMgsz8LTOzlgo4u7RFv0i5Z5vgwz
Fe/chKHxM3ladf2zKeKSBH2h+6qN9mplV15x2ENQsqQfCCDTkSOrNAde3jpaiLjotoFeu2CKW5Ox
XziebQj1cTfPeHaU+nbvobjELhy3GRWnVadjIFW/HabukJ3+DCF252LwnRfdpdfobRIj1ezcR/TN
59rQDtw9sDVDa9nOV1zPvT1VvgHsf7r80WU4dehZf64gARTIlk3KKahI/dl998KN7oKiBaEuMMsf
sgqMWm9IQXkmzAxpH+CkvDuwHp4TrH0fOHKvmEFMHD27k69x1zuFEmWsSi2MEGQ9CWCJWMM1trL4
DQZdG505Jo02ZTqKt/AcmfSZERdUx+VrFnvsp0U1oxtLeMDCQTeIFjscTPSEvCShRIumlWOubkg1
gN6HTmqct3s6Dhhxab+4ZDgSj79+XcuJnHy0FgYU0SuG+aBTycOti9xoxOpMbbxIx/aXaj+XR8nQ
Ef1I8wjp5VviySdCCc/Y0Zsvf17D5CXDGk8lkpytc8ATD7uFlYBjQaOQHyyUPnkGjeXlIaHZ9ewn
N9J7e5gP6aAgTRpfmNvHGet0WZgAVmqTT71rfgj252oNqdVebmKe5qgtF75oF4/bru+HTfiex7u3
ATLtBJM/pJn2jVHyd4gsL2JJMTxgIjDz0okABYGZXdh7K2vvc7rrG+iORt0c5/tFQS9tbTO0FAef
jF6/UXcp3HUrkPUgsKfsdW2IGy/z4bKzINnI10kUAq4lkM4RYKBifHhh1+Rbfg+JWwIbm/I9LXzE
NcIt7Qs0KORHDHDpVBncsLBrAkKjBPdP8cBK17iabIvdo8zJr16a9Fw5ZZKf4TW9zY7KjBgSH4zJ
5wYdxTTt+q9/cjOwhO5JiZtKhsR0Z48wMBZlICRDrKpjSfjfavVs3LzxFDXjX0Hco/RPVWAxcnwv
jWz0gbgqbeTbBjYuCENMXL5xO/+VjLXYuFndl2HniB8ja8qmSppPjXih7/CPKP1Atn6gqOWfwsLg
mHxcoN5VE60TkkTfH62Hxjzivfh2q8iF9Ma8gGN1Keuhh0g9YBXJLe0lCaSBgFTB5sYX9cRff6To
DItF1NoEt8oSP7C/p2/EJn7CqPdKdVyoFkn8zMl6R+MtnkEL4lhUU5db61UiH9RmFjJv9AJ0YV5/
Rrijm6Af6CJr6+M0m3/z6ddzjoBpXEqKvdWAey0MCmxVgLa8L/fmnWo3Mmn72T9eYl0cqgmfKb5R
EmFEjxOruGw5LxAmr1kHGXJTjKbEowtgfuYr5e8dYYenLbwVDdyXquKIoUQyNTrR/qtkjeC4z3U9
fkpNoVi4l+b4218OkQ15Y2ORDalDbaNvJb5fIeCXlQPSdKwCyV+GbqOroCH1014v2aOTwaiEn5ky
IPbnf2nK/Tk22S51/PZalnMH3cBTFSfXnoh5NDtj0+x1EoXvB8H0gD+Hrzpmxcg7nyYPRmgyZmxt
SIh88uuS84oQg5KyO1i/74TrcqxKwNxLyPLgcAX6Sxmx6PDx5pi/gB9gtA51voY2OHBlocCNdtZj
AUf+tRq8YNUkQXqoREpdkHmP4lBdMP9GGelx3u20qy/oUi5+K0SMwwdl//AGnmLtwxBV4750Suf5
PzPwmwc8CL+g7SiFV8shU7C/gl3ShcjCL+SjioxmRSS2FSdRQnfI3MNIzkfYpDyUSJqJHDlHGLWV
hTo7aYUL6E9wnDKzSn5uWdE9BTxXDG6wMoe9DegYqsBIdK9PHFSUgnvt8dVWVTqRKZe8THWl5bTZ
3kpJUV1nYmwSyF1QfdMmOmO7G3M5yHALB/TeuuS2EVfLw+c1LhY14jK37h4FbGHlfm6bkEUfTZoe
j24vlmkOsyopjuqUPItI648PUKQ4qbHOdPNh9jZyL60licSWK2GS94z13WVjFX7LeiH7ghZoNl9G
993RkgAQM+tVSGdDqQfAFqP2muN/4xYoQlYXLzrJDHXPqUMqOhQ0kiR28eCCnwC8eIeOXLXbfwyy
kHoGA3vYNrWLk4JJeL+yASEreF6MuMPopo+d2UhRCoVZWG1uE0YgMpdZQfNltfYqEherxyfez6+0
+Yo0b0In72GeqI6nMnzMCQ8gtD6bKTOvRekpQjaQ0cJ2pIWlz8s9wW8Xlcn+fZWMQokMow0k3blF
WsQWaQN9Mpp+O0Vxs3Ak3Mz+CKsq5R7745ySZ7q3fxtt/MlpCXc84jbnSqlpZOucBb9GfSMcvdRK
Cbp7HHWDDvIRqqqJRa59Er9It85D/qA+4hyBVRKfubRCgk3R5avrEPfPy+43Xh+b7jqOwZnV5RBJ
tM/BIO4taix3vsGskcXXUY3WBKTfeKgahJRb5pclJOvAQzCOkHUyDj+Ad3xGgvw0E7Dm0NV9HMqC
brxyFe8REuIXeUXaNsKI/GxE9cUmRvM0cQj19ohOnLMzEgIxzeKtLDfdTj86EfWHLDwJ6VPh3DQG
tZkXGj+QfMr8bmjXcIXCu9AzFU/noM7dlQ3mqpZdKdZIcBlZV9vI+dYj3KXKVXYZTwvWzj7eHC2a
xNggasY67nlDNklFWOLoYLRR9ygGlsZmEqs3rUbFxWSrC2t2hFroCe1IdSFjhqr95mtz+xyOMLTD
/izY8Xh/oQk0AVWcLncUQITnd381pEZzugEP6kkZBdfdxRzvO2Urn4vCuk2ZsU06GOs6Gxpc7gxb
DmY7vqh8WwLK/g7gcR+fmmndxvPGy6d9NnGrWEcFBNbrmEjv6hBcQNFiIsqMzsTtMmf+AbMWiy5l
b1yi/dNvVz5t1WXvuzQiF3fx+8AAM+MEP0/MpEJgir0hF/8iXc9A5UFQReaZf6WVjR9RNTG2r/2b
gGKmrr3Sv3JVDxgcp9UCW7oMBYAYX4FJaRFkFmJ2geoDMWBc+4W9q8aKnH5y95KPo5qmEqFism9z
c+wieTJiXzSaa976iisjGADw9f5uB59OrvDaqrvMPIW5ij76kbIiHeQvQ+H7n/LM0KxNpXhbzttm
vOKCTNPYSekd9i45VSfe4QuhsIalZXH/ZWWxNZAYSzOkK6oSBA8zS8I7JWbaxMpz+dx05qn4a+vz
yYfUPFswjkg0yGAczFO1ppCN9i2U7O1XPm3mO0bfXQaEVta8bOVvtu9fln1YyXpgiRkyMaE/cYDP
lJqwn2rsCaysF0BxCp56FsP+sRobDpIGEa+V+I5Y+NsF+oaBpaNCKsWGEboHuWEtUU9IKKzozRYg
6ddKxz6HNsYLMlK+vkoGpYrW+dHPyaCuUR036P7D22xAkq6nd0wa72XD34WQwlUawhWrWf7wnBjK
H9Zlyf1Z5Wms3ZCwDbFFKSefFrL8ZwUQPwDHYhTkjxJVovo8F7OhzMKdwpwvRd00sQfwRJpzOE+E
6vB1DtVdby8PdsZa/IeKWzNmDEWMBHhKTxYaWIOyXheQDohFe0Dt/q+sdHCYw6FbgSVbUgcsxvWp
U/k7ob++pPXIgkidt3nUkUZdrLlH/Gezr4HwPv36V4nHqzB9bT5ybCR5w2iqsE9Q0gTxvncsAcaE
LKMRLtLN4kXuNckRNItMDvt2n4OezPJBzM1nVfIrxG38QfPoNvVtvUj70+AUaH3LzME09R16PFU+
1kd6t9s/8fJKhD8uEqkwjQUM2Gr9/57i43Hxs0qEC5uARCbxcRcT3fxWAZrDTW/HX4gtTUnUqSKf
A64OukbQ8dDphoJVBESxbUIAxIIXdvEDFi+3aZdZLKpwcbYx0/rCy+U2LJJZVOQ7HFyqodAVWHvZ
O4OLsWVuTst9ZzutGHoYmPvaJ4tOnZcmf/PtdXn5yISCLF1o0SnbQHIPt+IX+5BRXDrFzDB/mWJu
dPMrhSyxVmdPPOH4vL/Cy/PGDXfxbYsk3TCF09gEs6gQp20wwCkXL9haisIhBMGg78P90HEcMK1g
ThVyf0CNzB7IRhgmELj17C3PS4vtBuxzLAjSuqS1FAbSc1eSCSryzm0+eesXYdHLNwwxw8YqwL87
lcHYZrlLP5hW6HswsdYrL/ZdJgl/MpdfZtkG6EDDx58pUwvHHnMTlrpq7PiOAl+9cHUyx7jMVWEn
+G41EB3mFZX68hoLB/1SuHszJyj+uh9IvLX1Ylc53vEWwWSw3k9NLusxoeH9e0KXHCYRbo8X+fJD
owXToajkctwav86hmKGXe2rQE85NQ0kqO2wm29d3bR/EIatkGxfDdEqTYNU81wVqzBqOHvnah0Yq
jLQLPLXhffY5kpSTYcfPnRsKuN7E32sE+w/wrmpX+c8/LQHD4pW5KehCLGQjjTxF/McFCWM/mqOy
99J5kIFN0fHo92kqla/2MF7uSDuLE6JIb+QVbDRq6JijNTAWrikUQia6G+dc60PadzMWzeNMY+bv
YjABo/Ck01fHSbOFbV9eVUaZ+304sSoSuHD3/vFB1wzXNzVb8mSi/zZIpQw4/9e9/36ACteUT/PG
R2TkTmjdB/MHJ6Wm768pKJZ5b1TyBa1J2Y7k2itOo0SjUfENOcSoya0K9Gj70S/W6T23vIJbn6tE
cXkaiPfy72cv+YikwPV8wZI1zEXidvrG3vfZryiAAp/WPE4X1Ot0lru6hPh+WTBLFG0QMGPcSzR3
1X4ypBDyUPRHzuZw6xVteOpYhrhFcVeL65z/wGm5fROrWCXl3VCRFJQLccHXjSUlqj6fqLJPMa7P
AsZEbrJ2ArCE5t8PPNN0pQbGOHD4iduw+5ym804cZX/bFarqWjiAOAoqYyBc8qcT+zHSMlI2RLo/
MIkNAzdKFypAe8S/H3oD97rPDtJ+/kvqqRuxEeF3llWis5jMQogD4sd6pR8gEAGN/8ov84dBgn/W
w1gqoRU1TjuKspSsOg0dP6F3hxZ+zSP9Du8al8TKQiH1vDa/XzPWBdjrmR61qqUXMbHuY//vKzeU
g2+RtcFlU/oK51uaB15J0746vdTGiT+RT86oBZoIZBG/KWQru5rxRYFELTdoP3dtzIfcuhBwS0vq
BiNPdTj7Ssre4UEaw/JNz1wE61G/nt9+z4/hF2yO6uuouE2twFrmdT1ykDkmhD8FyHpeQ055ploX
26Qf2Rbq2OsWszJxFgmtZA23B1V++Ypl7ozuOhU5RWdE5AgytuPE9xfro/40rOz7HxRV17V1bONE
GqZmNrNFICjAnBmTZwkBevrBz+LBMFKfGr0UO4DCc/AjOpd8Zk00ZJzAeIutE1smH9DpdBUFG6M/
Po1hqSRNfELGkiJxd+orvcjsrFrooxUkzsGeQvBnI5hv3ZXIRR8JHLlwKpFq+PX8aHAMUovEsVbm
bGwBJEb2Yg2WfFX6zTVR0VZkJhwpGMnIgJjkju1oe++laD6C9NVuOp9MMUa4+gHl/o7JgD6Vv+9/
/Xy2hiriXEdAGM79XiHU1hsNnZVToga4XPycs67zA03mAnoNwHkJevMbBSNN4KbyFIJKXVaUz+KB
elh320+zUEsCChjkAEqr8fX2XsXl5WGsDfxoqwXEUbXhRf+EsM39LAgNjDpkac7AGcaVSrJ4gdtX
gT6/Xz4UmPLLtXeZ/VA8dTh6S/XzWVFnimc5i5yoV0BKTff2yMX6jfI+9+PSZupPjbPLfLxGuMQb
ga8fB2dUVQrjiaX/tGs0LKY2M1gA7E0ftO4fCBPf+ANe3ZNj4UGhEBUsLvZgn937K9bNab/DFexV
U0nzn9S0q3zgMmgcmpcbqHGjWDO7dqQ0HNtJzJ2KlNMLVz4J2Zdqd13DuHstiiYTSKn209BlQiom
j7Vn2N/Pex8gGYYjGVld67NsGvsyr4jQgfc9B3gQrjUVHoXcDHrvTcP7UV44cHNG+ZLzEfAHAI0/
55EH8XbyXyG+MTvN7mbzGXqzHcfGcA1kqH/81UX4oxQPS8V/jTQ0hOJIfPVyUWxtm/iBF17GLicB
mt7I5l+INjUSjA7u5RjkQevPFO2Ob5IPkrZOqDSnlud+PNZySoekIKVq1AZ5vSjoLOlbp72rib0u
9L98BaxOgY5FbF7P5oVFIwycROFQE19E5AFugYBOWJewx7bAieLJGX7M2T2TolWZ/qih1u29iK0/
sEtiTrlA6Aot/4+uzSn1G5DfyTwkRkDRzKi1JEKVUK3DrrMq8+7yJpnYklAbCrSH7xpsFzIl+l9W
jX6CMGAV7W2dLca5mWf/aOr87u5wXoAeyR7XS0/nFx3mZ4vhqrfJyHOrh1Ib98kSRRbS1Jl55Wba
70lsCxZxOAevMr1yd5KVsM05/Y3nBt57psLMsj0ZgFNWY1bfArCSH2iRduRJCIiw49mziN/Hogid
F+d31tw9n02cJT66lLEJL3T36iROxkUyejUmzn+ml7Pq8TULqqP7VINPr4DO2m0SBwXsqPQOnnqt
Fa8jJZf9GR0rWRn4xN2Gm9dJsGj3DkT/K9mCMZdxbO4SVwx0FXTBdcNftTK7/JhofOhWFJIzZwcV
XTj+FOKCOfk6wbWpDk73nNL8PgUbGNuwQRL7ZsQvnSgFUKmcq8/u//t0484nqQsaPouLB7Z2H5tn
tLmEGIlDdhNfJY8Dt46MPCpINVD/D9isJj0YIF1y4igMFsPmva78FY2QsjCORihWvk5xYRoqhzjh
ACPhOnRRBd3p9vsddPTJqEdTDO13vvKfmuEFuqLMRVGsGefORAaNwwtzffaJpwMt0HuTqRqRkpux
aOhIaATCvdaaCvTuU1gTcuMLln+wZ/nfLYJ/090lRLciQ4F8HiB1dJYA6TTciuqgsypt4X6B/s01
OrniH57g4AGi8IpXsMGNdgnSJg2lwS8XJpvVFO+h3a6JoAN55dvmiVCaZ/NyIVkxx5lz4wqN7jpV
tN5mYeD36oj/WXQB3V29WN26ELrdxxxRU6TjFraGCZMQ2h16IWaRwCu2ek5icF4VbBdbUkBsCByt
wThEUaHh7ASvMFWfbpdVfi1oGiVR20pcNKeUYgXkxhFAhUuV991gVRpGFpOyNPrSr2mel9dSzxUf
IqkAB8dmkooJaQNUIWrUeVYnDuq4/gEMk8OYwP6h68zbx991GGQelnL09+v1uAYs0OY2Tgg+Ppiq
hBvBEP0wlGsdJbWeVpX14mfYWjmEakj3YdNc4SrDRk4BmPPs8kx9iRlgujRdfYCBuNvMk1enR1P3
BGwCen5Xy5z56l+xqgPbf2UvtJsNyJHGzjo6o6EMaN51CAMr+3SFA7srmTfg5FxIHKnB9eQ1HTv7
22cmk+nHVjXwAghkuyuLw0/BE11SDk/Hd3G6WEWK9MslNOmLg3BMCvZ3a/9iD+y+PPAbPHrl8n1t
RA3BrvSFfQL7c3V34nm2d8FIebWPGXGg0JwRJ+K9KyJsyd+b0qqh08+tbGzF1iFV1WpEhJzyYXko
GOzQH5+FChMOJy2303hlMW4RljkxU2VixIc2WJ62/B7jMILM4rsmXGenXO3QiW4RTNCduBcB2MDP
mne6naSg0S9DI7tCBguAKG4gouwUFKlF8S3yY0YmthEKl9XraezllDLFoGDCm8qgD+xh6YVYDpCJ
FdVWTLzus7Mi/MgCOakBw7rM5g22q7+9A+n6rc3fS9LA6k8tI+/36izA/HF4drYXqKu3Bdzs+nRM
/QceEyzoaCeUxAqq1ufWN1F8hMi/sdQSAun56NUhaNLVvtEB1nhba/PbZSmpVjZBKEwnKM1xXj15
EIzEawHU4oyJz7f8O7PTIDaIBNDmLWFwuAAfo1RsNSqU8AHdNj6RC2IJiqZfAfQ8eriQxotajG8Y
xdMO53Ws29Q/H97gKAkMNmv02LYR2EDbaB/phk/eLMALZHkA7M9bWb87IKUItGBvFIibw9WdiFAE
KcWIVdSNljl1H30Ost+QsuPepsD+bbEeWKg1Ici6waGXnmhEd7RQThwg//kPc+AFgUb0SKxggdB3
lOPKJtrxX7IQrTGMeewKuZWwX4r2jdUAzbirV5fFLEbL2yaxirXp8iZm4sTqxpaSe1RLWowDOv8b
A9dKV0XAKrbrpxJcGhtp7r5BnTt6tuCE5MA6eZ2mbCAt7IgMZZhUT806+AEWpc6zZTRc+odhuJtV
v8b3O3C8gN9MpkNfFH0Fnwrt7LIwvXaV8wDp0BxvOBJEgUuvG5ChaPjJo2DHDSIbAY2XQhdx9db9
KQNw6mk0ok5RyVzVZyujMqxTUOuEDZmHcQW1JVzskYeQ7cKce79zH6Jm88dDtQlra9+y9pG9ydn2
nG9I6cP3uS9bdfXBa0NoL+62uEwgy/KojbFznCuZKOqQ5KqtK6Wcu3h8DvpO3XTH+VTMC3dQkWJp
Ojq7dcNLOZGPX+xI53H7ZS0R4FbkNSWC9JKJBAKNvKB9VXiDZCLHTrTkXz+mJLJFSFC/MCWw2XxD
hj5PQilJmqVtdNjVyBX+hoTl2p3pBUJmOLo9gdg+UgdAQdddIzGQ8umn57QkOY+qmKZJFhlH9QNN
EKRzTxWdWwpqEhxV/zEngF4RjNSm8Rl1bAKEByEA7hsVcnPc4KqnMy/Kj9nBK4N56mdafK/WBNP2
9hON1u6oraacUOzkrMy90dP2V1qW4gwxl4ps6Q4mqtaMp/0c0LzprV0oavsgexIt4DKwezbB0Ysv
rpH590IJX3ddGvUlqBLU9LpwfuTdBfjjmELIJLIuboNtTfICHcLZkEk5u8lsA5gG4HnRgyKviPbX
SQBBkx0+Rt30pxsjJx54Tlr67QcggVZWNNw4jCiQ98X4TdQDfNyikmt1z/tUikDIyT2pFa4xrTA8
88GvS0wM39YliTdWORvkzyIoI8VpBB3lngOkDLXNBIKUw7S4ObxdN74Us0THSSr1tltGS+otlHZq
HbGHvlBQDTZbG7t7eo/MEkGdI3eKQDSwhFnQ+Lcg1/eWFmOsyIBAudbgxMMbgb8x3F/mCYNuOBBr
llCXRXq1hsfYO4NPN73/ZZTBYL2JR4KTEfleDe5l9hibUDa+DJUAhi6yJ/49cZCK9wL9UwfX50k+
hei51VSxJAX9LZGZCihbus8Ejc9fUw7C0CRY48EWu/TS+X/jgFwHn5FlgcoIwnM2NFp7gow6tmQu
QQiFBH1/WWTjnXaBcdASCU3oVAgwSUYvc7Ivge3htDbP8fHBktBgZITTaAFtFpR27Bofw0ws4SQ8
0RnptGj3u+UJkwUgBtQF0PZM3+7XPNGQGZhVKz2qZUdMbHPfcQW6U0Mbh0TCoX3kCjEZH5Jo7LOB
Qs5S9Zx0w5PwPXLzjza+P6trb2krYPa7Um4sNki8D4iYXJtVxtkt/0J11mE3BcWzseI/cZLZb554
MO0lc3XWgEWS1rv1Y6Wn/cDJMlAlK+pnMZxZZz/uasoapao6gK4QvBiNSATwkID2wSOTs4cupwPp
gg8p5jXOZd7d1kVis0gwZqaV4yw409+C9F7tV6LgTB/OxbbEqeFe4lAZt8Czm8w4MMU+IlOvKZ+9
FW/+wFBkqbU1L7V4+z93jAYkOmAHY9+wW7WvM/bpyVaeQ+sjuvvJ5BZzNz0k0oMgFnH+1IoA73hq
/gfJCtXD8nrNujqylOQAg+/OmbPeQhlZ9NXl2Hr7zDor8fKl2lYLr05kfPtdIodAdHipjhr/B7wj
W9sOncixkxIGE/eJPxg+IlutndOz05krqjL6rdTDgNFOL2eK18Us4XgrJaILdsxW7rEi6K1OO6oU
8zpqZV5kPHtvt/321ctp/aaEsUYwqFJ6xAZXMmG1aBev/0P0sGD0qZh7UGrc1uFxtR4hIvNm64/0
/aJ0N00EdbcpTupPDlvPT2jd3hvJNEuMsYiNpn87IEFbHuHhszlbjv2GXu7pytLPb752+IAdW4tB
9dPQJOy+y2+tAmiF3Qqd8XbhwbcX3sSzdaHRmEnwDgwYnzOB1sM+8Mvtb8gaHr3gEC/n8ZZyyEr/
1YuFm6bV2SSsr2/xwaFGQJRpQPchTXDmHlcqV/0UF6Ip8D3zBSxQ9Kr0EzDDdqC/EWiEqtzGcYqR
gOd1qiGrlX9qcrru3uroHklvnAm29ko8HC38zU69SvN3aYyWsTgpS7633zTmfIexs6TPv6K9hq3d
GgW3Wp9r6VW30p9a7dSpwYnLzfyl7iM0Xm7hxz7YxbdrTc/YN5SYKzrwuZfHSsh10i3uHKbFKq1L
SH3IcsOYU9hArmnp6GU/0eqHDCiRjbyTkpBUaikZDwAOsnvwO9eU4tcf/gwAXGGRHcnhdoFFCUzK
AHDBvtoZ5GTIiB8mALKrk3xM4iglxeUCs9SdEv++QLV3xscNkXx2j+rnIunjxJIdeivRVT/ZcfW1
tcRVULXipQCy80A6l6n4PJilxjLGEYt10WXbFKwxBiiwm+jAaELKBDUy8tcRIS9lLgr4QlLj//C9
rRu67nPXzPjegmZzUXyRPXVRnkbCRIdBmKf9UAMLnYlgc5rB9m0hpRwYpoVPNBr0pfDM8QSdnaLZ
ObCzVi8t3HeImpzUTVGLB9pzDf22+8+6cQt/u0hdOx+0hT7o609iitWMR7jpAwEiJdr/JojsR7cV
2gWnQOGizatAoPg1wRqBFkOjTvB5DJd/XbVfYF3kQzrNBaF/ZuAUyf8uKLLQiPpILL45aM9ST5yz
lEYuA5278uDqWC9AlGBSKMZhPLyhoEa0Gx93TJS5jGD1FDWlWru243vTYsoKAx8WlRhSk6OVF80Y
OYRgdlaaNHeMVjazaN2YyJ7PmRkQrGEH6NONoTTYGtESL3wEa7MzKRjZdADmuqGBrlMNgthZEy1I
OAbyGN5waS2ySIx+k8RDbdPzjWdvLBPqgDMiFfBLGhPi4NusX0DnrQzvLJfYQRPPKcMiQmHnTZnR
ZzjT7mIMk108F7zCJ3XCPYuDczB9pAvJ2nlQDOv3jSQbnhSFfPGp6aCyB4VbvHH3MbG0kO69vggV
z9d/LlqZPdhOaV5xm6nI+qAj9Wk0PDye2Lju9EVYnG4/afqhZOjdNDG5YyFCPVRCPebhjrpZIyHb
evrrDbYX0nh91g9ScXU6Lmo7sgi/kOGhb3ZvWFxt0Kes2u1OaF4pG0Xa4ufHWMn/NjQKYn0h/UFn
g4Q/EWf9gecR0ds3YgPZPWSgBVHPt28pLLHs9XGyWkkD/aZ8fGmBo/zWlMVRq8Va4uP6ikol5vMB
q5t3Y0ZWVBbcDbQ1X9f3pjcBfZd1O1yPs7TAZHCZs6Gtsd/waKXVDN38Lv/vK7L/cdD5oT+iDEUN
GcyqB60ZGmrCSsuqtupX8Wchzer9dc5VeXSH4HlTxheSC9Upntns6eDy65U7g/iUgQkBQZ5r3IPe
iSUdjhEJWorw2DdD1ySWGEJfTKoKTHZfILEVZLRyL+/wC171u+lYqGGVtTFTRvIZjtuN09NsiXjW
2ebzJjOb+bvNm5tJY9+K2rKRyqcd805OfKC+PX43br/jD1LMIDfkjAmBbhbvRNm5X1sCl6z6TiZN
JripxwscO4kOMv5w7VUJNtMEzEr4vrkBh8SNvD373seX+KcZrtWIzaADowJ56IdHow839lEQmdaG
H/dwaKPaO1gzHBsO49SWdGQEXBB+cEL17LF8hc+/03W5Sjacl10StgMjSSkf006bcMjG7mn8wqQq
rKYoYCqzSreP08hk0tcwbb5BgBq4V+DkhzTRozITNqL5YTlSmsNHZnbIGH13QHDyGKUZxz3bCFrx
CurMkN+0akUzyrwcljniSlfBVTVAGtfpSfISHFB0ZuFUftjXBXsxo3//9uJ4+inoMiR8xagkbuUd
wafnvNadInlIt2xWB5QGmL6ankWXsVGtFcaRa4XCMAdlegB+cuiICQfVMKwq7BgV0/URNtSRaINS
1baHY4qw3hke+tL6tNIbljuhfnm2Ky/u5hQhjlYlq4dXh87hd3BhK5W895WvLv3J/JB+uUwzEhAy
ZYHtrJDFjPxJkP7n5yFsUonsnGeylqOlLKKQ5LQMXBhiaQDY9JAFo6EN+LfWtrmFliWU4Ce09+jb
hvkmIEJYXTq+mxhFpNj0hs/Kt2hgF2ec+Po5gyQQcq6SGDzfwzSWt71E/uauK320T3jhKATr9RJj
FMx2bFQrq8Ghr8858gtAKBPBssmhn9o6eksey/KaqNfXEAIUhehlc6TqKs8DS/7gQOIbuJ6Bek8Z
CQqYG5+oF+qs7YzmAvxvKM1od+k/0TQ0bH0+516TBC0r5eovPZsf4+gZYdWUxI3CYMn3Rev/fPfb
Nlcn2ToSCUQuom+IM4gEvP8CAcz1R0AnzKORgJBSLQlUzgdEpmmQX4ux+zJCrxF6bLD3fMzcynbl
41xr2mSStjZ18joV7Caj3T2+BbFXV+zo0oYyeoSrDVACTVC6485aVjxY87Uyp8f3sTnuf42a19XQ
/UwMF7DyK8HvThwpHVoJ6NNNYahfP2aR844DR3oZzngedlnT55bzcm7witXGK6mOx7Dmp+PFazNk
GhIuF2N/K0JZEoQIyt9VV/1oEkaoIwb4RhGX0HDwycrJfLqr6EN5vEEkYIQU7qixnluJbS8dwCg4
EMAUVUOsT1//f6wuBgI+B7Gkpca+KYotmrPHurtqRfjFpptUqQkNVTQiInX4mjhfypn6FOIAEAYY
+B/4TLyHeMzFF2fh4MGj3K6P8I2DVJ4QdkomC5HnQqDxyYG0aiZzvOI0ld/nJXgK0MloZ00yMSWy
Rp1Bcd3fptkiJo4s94F80M7B3bT4X5saW+9qx8ed4ZEC/lk+ej4Owk/dWJEcYWbBg3bEUeNT0Tep
dxIYsdaGCrKbShJLcyyJbR8CBXjKgeNrGZ8rBexg/TEKid0DXnyfTWboZR8QpU2lvOUUUqmmCc4Q
oUh1PiWdE7mDANtrEZeM6Ylr1xGv+V9xhMi3Mas10R7ZywwExkfDE8549xCkEKpHni7xLCx9XTae
8uc+weAQ/2ROkTIX+pH1IJORLucX4sqdIZ8f19VLe4fHqOwXhD/aPkVIhTStqtd5UIRDgJI0MH0G
DQI1plzOieIZ6/0MbdZRpEiHnzkQzYue2D1IqPwAU2FFroxAHxHuK/o7hNz4TqnYKgWB+DRYQ/eo
b43OkEYwT4Zu4PUJE42138XvFCawIKIE5xrv161LxG4dWCdBx1Xp+6UwJkXA4QQDJXGJDlN+L5t0
ju/OC33sHyT+ZKzbzhmOWy8Bj5pQL2H4dg8G/IIXAHMCiE9ya/yxbAg7S9qk3+ScBm9C5HcaciVB
8NLU+sFhqLP2F6LiPOWYhIAJqHxTPeuFcpRaI4K6ZfBCEKCdueb1YRY3JbFGxTFXG+VeVMtkKMN8
TZ2io0I35+id0od/nygM0ly/2YTUA3BempkRgTMm512hJuXUaFBFfnYK0QQkRfXXQh99l+ri+k+n
WGz14/uyILMsgIDh9Ll9T4rk/pn7YfzCVuHrirdKxVG2fi5QRMq25tXITF8RAdOwvT2+vx6gMvWJ
qnGfnIf6YS1szancaZWr8fTYoZE+DxQ1X+zPfMhQOTlPSUQ5ZDWgvxUNbO7ZmyBEMSVdvYQM4VkG
2behcndQ7rezdpajVpESRgf83+NeVveaZOcwEVYlYDnuouawPqbplFt4w85AgkGbANvZjf5VFC4E
pjqGbxS4Qmcgt9nTr5kRPR8TZYCb59kgE5W3vjRcopxSs5xW4B9oGnv4RrVg2CoYk8HPRJ9mtzRT
Nut4ksN/hO7IGvxqXqOvZ3jBaOjyQ85c9wzVVlCqTALNnVNkh6yp9AFWaiD71L+X4Mz2CGXZ32jE
JlMJ1Y/iHWbAAqhOy5PrwRGD3CYq7l+wX1fky9rMlpzIVjN6Z+11wPGxcPQ7mdoDUwL7DeY3AFov
X3yVsYea9QMnm25MWDfRALSxqd5iv6+YGjNHuMArWDzt1xZ6qPHcLPKtueyH8LkAhb+PEpAOTwMy
jaStgr5tyujzaPKZJ5ppJqEFxYNgXjcAkS9nm5skjwrmiOFC4V+UAl2dA9y0Oj8djurfSX9Wa3so
muj13SfHN79Y2tjzUcHEl3EiK1Cr3TyDMzFkU+XxZ/owm8CHbjmb/enBf9IXQsdp7+7RqO5g17Jx
hjRZvcBDvVDMhq4u892RuLGSYbSyDYbA0H5wSLkacl14GQ4yTsgFFhrfmuyK6VFw45/U4yLhIAXB
Sau60Ce2YdpqTY1zv5jRT/+EtDPGlQ4GOtQWnCXjzXuD4OeYGRRvvpRViK2bfRbza5+CYs0lFoci
Ii1t9qYJjxWdCosShoWJA1b2r7xTbHfFTu2EAs9XgeYw6wOzgGlo+x0nEvJuWxtzDL5m2GzJrCpk
XTa4XN+rKDmrheiJIw3sN1HLqBVYmU0P8NansCZviblPmBqCXz06T2WHWqNHIewcMfMNhHCUNChQ
/a1HYKWY/EMOY4yz5KQFzk18fSbSqhZ4DaS4HjQf5pnuyWuxrGrY1RYQ+XTUY+1B5LdG4njvGygx
tH4tHcnLQAe9641HBfWYKVjeGjBtIn19rnXWxWD41nSEQCTemYAc8Mg3iY7gFI8PY4zqaGCFtCMs
YH/iCl+Y59+kGvqDrCagSYPCs/bkkmvOHhEp+IANz8BS8Ty8lgvPvbL+qSIzpyClH+si4pKPMsji
+xpBGvj0dGZn1jRl+ZjEyOxATaGlr52mSKkTK/mVq/G1TaIAJgyqiQac9fYlbPCRO1NY2ctwTBXd
l4nYpn5BvmM41HeDWVb9fybnuaFM6jdb5wNlPLHLqMbJfLgPrTdamaBhyqNdBqMIV4iKwSmZwRjO
FdcMGJwZ+yWhGZUjIYewbwbUytqp2kzt2cMPLULJwl1Gp+VXeed0bajLYD9Btredg51PPA6YD3hO
NLj9v92+jnJ8IqxMfnnCxSYjg1oWRVK2U3wxLqv/LCIwn/TLDsjOY4Z+KqXW0Y885RNRJ6lLLSq+
OP/4A3/v+8kT+aPXPHv37mTbg8drTcAqTiUYJytN49RC0JmaWSCV9kQMf1HMWJVlABU5Ps+Tkl/K
434BAqm2s2z+4O9cpilxB8v/dCf0XKTA2rBRIJ9W7n1VvW0hOW2NWZuzIoaCyuzfIPwwOrN5SCXy
cafYABQdFxCF9MYpEx9m4MTpN97sJdu1Mo0aC5FVwTVlaWuW1RAMarWsBpkcTg1BYKTLkBv8e8vF
MlNg5vUuYOQ2TBo1VxpFw12wbN/kLheG/iGx3totmvM1MuemIJw9JjkMM+LEBW7bmMnynEkVsXFh
CwX99rbFtseyZClYK7SEurst5k/P6Kw1wYRNkHf7Kc+AQ+GzAL92lJ0UhaBrbCI/I+JXayfquhWe
9sy6KCyYtjbsRU6+sFH1Kd4rkZD8LS97qeeOahZXMVlvf/JbBQXGV/CUQ3aW98Xbd8x/gUyuUaar
ayn+RCjo07mf5qODjMFE9+k9H4Lw2LOtwq1fMfoZV4jFgqazL+kCLoKajnJEfJ7G/+nOySMby5wC
y3QJlpi+sEIKuz25oUyrBFnuaoXBz7RnCn39+eKj2K5HKZVqR+kAERjbkyH5shPCnoppfDTyRPWI
WBqLLKEvwjvnUMEG/zw0T/OxJuc8PYrLNBS0mgcG2r3QjRH86bO5Imn8VrbtIHTD1n67nSAPaJu+
gW39vy2IlgivKF9hd0C/GySeeaeBevO/gbLCf63KZlRwPy8WKRFQ1gyns5TTw9y6WDiEAAogdb+f
nG5Yq0Sskh8jcYrp7iHzXKSS0DIM1l1bq8emblbIBxCSxLBWIEofnbwZbSD/guGwP+nbwVutKj/P
l1pAo94yp3/dp7oDQY1/tsT+I9RXsYzBHHHlz2IgBsabAqP98W415RhHvn5oBZI+k0mQJcH73yOz
HQpO+Kruoa7oF6kQgYlZbLYleEni6b9tfGjx6HmwzIoX2GD+HuQ2cPh8M90h9PTFouvYcs0bHWEs
eOZsrsi3AXxRGpRfisHx/7bn3yjyeiG+6Bn3Ib5PPtXyS674COgRAf/NpLB2nBOKHPM7q6fSPBNa
7i//EYVTTeJTvVTZHkdWguZrYNaDEkEc5ocuwdlV/QewRhhBrBL4k6E6p60TbCy7JDOn96XKrNYi
l5qBqLy3PESGZIqkr4ACFnbITT6nGFfUzt7ZUyn2016tBoRYD1G6trqgZ2JQQVpOx83hgvsQk9rx
1/S89iXrA8VpVtGuOPiUApuL4LkmJd+3VoV5aSkW+SnMwBzlZ5uYlWzpXLHS73J0J6no1MW7wSZi
E6IzlAqgLbGQo3cr3j3AJWNOT0sZ0Ia5qck6QzqQROnrXlhUnAXTdggkQ6ispjSJx/g0Iigly2S6
MRm3pN36YG14ZZsLTWnsETGvkdJM75QGWcrqX0w3i0EUP15ltJnNuCOnv2Sqohd0cm9S9TH0cbNJ
IT+bXi4cI3sT+q2fmxl4fVas1FOI4n0aSshFbq/DIQKQ7leN/nmpfYi/miDRfscppMGHCHphG1Al
APJH3kSO73z4EYimQDPqbIj2vCmaN9lJGyVJTkUcg1IMgqMo1pOduMBYVkF6/uZV6xqwCT/MWnH/
C7Dxq8vqZ5rkjuwD0PRAqOoDuGE2LUS+y+JH6M4AiQp4mNkXU80fUq8ycIul6dKpfD8hM+EJ96Aj
LE8ypgQgAs+N6ul5ND+guAhuEhwxJdVKiItEEZ/ImURdhuu/y8TUBQl2x5k1zzw2XgIReb4YD0+a
bnoexTJN7B5W3a67MVuHBQbeo6cnT0ZRtRBlpsOJGPcG0w71NRmZlK02VneEgezxzY+BpMId79FB
3jNViulNOEL1EWqynGa1VZH/ozB2ETNpcFERly/v9B+P7LC/ENrUvtrdXmWwXFP3HRodoUiSlVRc
UWSual2ITH6lnFAKwVTslcVIDMqG9WvRFFl/WaA3549wDyiDYY87hoO1KGFL5QwflqeuixlZcUAO
PY93J2GG3nHVGUHqDEb6vDoRj4o/oeO4mK5yACjNdgoONxXLULA/Ks8CUOJALv/SSSpa9rjCNade
/ArEwrsca8K2W106FHtZ14rw6HpGBmgquDEevEL9MjEOW3Pc+LLX/WDjuDeesItoZAPDVBkxRBaz
0Of9DdtFURNO1GKuQFiJ6F7pxYIZJfSoRWDx9EYnUszK37HO+tJjjW2O3RdfXYttqs7w06aPNfEh
fnYMYIPF6F34EwY8k80K2/CVGP4IKPkN9Ogc5VobvLa1HKFlb+K234XowhSHojPIQkbS5za5iHps
zp0QGsb2KV8wstWIVuRwATNbfiliHuacSOB6A99WhBKvNfRQTLFnLHE33Fik83rjy+1bQal1bLug
wbWix6BODLG9Mi5PwA9FEGidEpT2+HfdSUFzY4wa5XFSyr8/Speh9PHdVYOiB7r0oyqOXfoYD5Xk
75wX/lcK2Ysca0jjoTTWgkDNmCFjGFMNuId/2vRPXQS2K3KxXnklezNye2Cpa0pupKrLn6XMowIj
7euVCxB08tzy1/jU8KlmB/FRWkMDxhrvinJg6lJ72QeWA8MerzVCAZWUnwBDGLHSEAbon36c6eUI
cBAGi88HSmliOyx2T8G27n52cXJM8L4M+rpLBPhoO2ISv6aldcBPpZvD+e8ICmo6gLK6GQuGDPAh
pjFrra1l2QDtIqzQuL+00NMxp6kCFmWHRECiI80lcIey76tat85L3i/maP/zlRIni3s4Z5yXkArn
KNmr/g+k2HdjnjIsfcDvJoxh8qclyEoTNsz5Q4din/XWY7mQ4lzq4DNp37hS0I3/oCAT/G8jS7XD
8tpIqh+ltYL3nGD5lDmQxn9G4BkBjcbyVWHHDIwnA8tKV9llDdIM5LfgKx90DDxXWgheOa4j/vsS
5O3LuYcFTcWWisXBBeWxJ/OEy9SkQKLvCha1L7ARu2qxTFBE8I6z3MyAw+CcDeR4lhwGQQdqx6/q
19m3l5/FzwbxgikeJsxF7RPG1JGpXkTqKHCfJ+g5sBKtkp0AqDA9Qjh1iixfUWYrbE4oEGr9p2l1
U0w9mjQYDDgxoDorsqhhVL+rGZ9UbXLZJdmhK78logkXQYB7iNQlLxMOQsor2h8sbV7N1svo7AmK
oC/OfHb+UBaNIIxskQ+92kZT+EReDjfQH3TV37ZejPyLq01BWwAtDu8zW/BAR0zIQ9u7JXXpiT0x
i9OTBm6n484bcvfdpyJNomT55PVirnsLcj11qP08tAMezyxLd9jSWUm4Wt0g5dXYxfJjsBwhvBaJ
vADw6mfF6/djL5YB+4FOpb4SDAR8gSCK/ZT/JqCMNJ5iMQ2W96qm3Ju4jgneDGsaMiGQNeJy6/nw
lL2gBXd3/nhImqSBkFwHCeP5Ftnm5poqyyt11Uo8YEMKhNvO4IhaFppsdPUJsXwI1YlJVHx7Ffwx
yag5oaYkRo68rkJ71vBrMVajy3xNbng/Om4o1sYrX3CLyywe/6Yfsk0ldDRi/WcSEkztn9WH/KDn
MSVWW3e97wfGvoGyXEUJwQuAB8F7H2iktuzZ45dCHdnTNSYi7oAykow0VkSXxPeASCcnaxe4eozG
mqQVf7MvM/P+8dXK+XGz9dWpnx2xnD3wxltNe2WizAChm15ay3EEyQ12x8mbOOWZV7BcoJPrHjzE
dApllsrnglXSYOQ3UyvGA7q+lhfm3SZ6NJ3VwyeymEAfaroPzR+nEsutlO/CtkVwg/DIx/hHPvf+
jPXiBf5j43yUUIWtgubqYLN5nAvNEhnQ9ZJ6LWOd7JnGc98dQfH0G4RUfG96wbZsICOVi5dkzQnS
QqHtzad9UDIvEmgu6E3BL5NZfCqnawjseBC34Nwo2GO2lH4mokzk4HdjxFf6AOqb4qy5YLmu4oGs
M3a5hE/qSB8tRa9tp+x8Pd8flz9FJXVDp+awSILM4uWWKvRXt/vDGJC7czzlhFBeMPU6B460yDZO
TBunqZj1aenIOtaBh7+0XiT5frJF1ZA+vyjphoGXqiE4258nVskwD/edicyn4GRt1ETaLlEMhFhl
JWxCj+t0sF014o0dU3r0EHbYBTksxsP40vvwqJHzsGt04QemKqBb0g39Fp21JsY/j1tGnlzhxiWU
+9d25Nyp+TsupolLLCeQo7CQ3s+022P/6yMWmiXUzaxEM1+1VgTCfzih3RlanDx2cSwoSNJyQTnW
goZEZ9bAQ4EWGnDB/1QhcT+RQrnEQcYh0Av1VXr2hUo8FQYIdijiQGhSIYzbfZ95f2srRgzuNSt5
/FqSF9NAfU2AsxKF3sspnCndUSqNe9rYpf1TDaEmP80MqGOhkeCm5O4dxvtPzhd26M3qFDLIeLUL
GGZCFEdHLTrm
`protect end_protected
