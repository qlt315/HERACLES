`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hgCV5/9RQ4L1ipYLo+sQc1RT1Aj94sjqVAuLh0ATN3WwNppunIqoKsxsijfb+RiFa1+6EkSc8SJU
uO4vv4Meew==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rsbfm2Fh57xF5VXWUxqu9mFAkX+V3TAR7PT8gZvQDPftvBh+mWLyo3WwGtnn1sIKov7pOeSevB3r
nirnytdvFz4UkWYxbK9m3eRNEWKe8ldtX6mLrTk7mXTqd9gGVl/SoBWWjRBabeJ/87U8u8BvSJBr
eFXJrNJwOklNZVRjE14=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZaOlUgItZBccBWJnBw+RAFrFWp0TcfLeVFCV0yyIAXJpvsBWtvc+/sEsO9FafqJDliWjJQq048k9
mCONVG/0y2HRrK75BR6YrEt/CLmeOpkIXPNtoLjmfGWKqmz37iOaHaB7Pnv3FHubZqeXnS4HLoZd
bpWZsjxBBCOafZTy12nsfWDErKncYPnuXK8aFK5YCqvsv/YyXGbs1benVqrriUbzS+uV6bl3hx6Z
mk1ky2moo4+Y4SKa7RlNQqyo1znRKTqc4iVJHcLVQvs5woHlUGfcxq3Esxsb8ip2Nn8z4Jgy6xZP
yS1gA8GbOfyzhuy7IDyyIcV7dD10JQ4EgFXmuQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b0L1m0tEfkDx7jSmzHH8pz7ylu5Wq6dftvh9InvtaKa5eozoa/EcOJa7OLuyW5q8Z5ORdB5UbCZ5
WohHSiKYkXgL7JmBiXmH4Aj34zp2on23oJ7tbjd/Q3bidDg45IC99RirB8v/rQvlyGtUg5cnjIQO
RLs/Lbxo9bb10IqEMVZIGTLZT7y0ORIqit9e8fDEz//G25qu8WE8oD1FB50Jy8n4HUnotcIv6gWY
UfQ77L+FFja2OiA6wRVH+8ykMD5r7GoNNM4i9IlzwNne/x7zr6NXvzfvPTfn6YBDT0XFBbbtaT0n
XOJbEyZeLV9NOxWadSD5KxskdYkBZ1pHhEVKyg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YuFiAvlO21jQ6RHHHkclDke0uAOfGpDfTIq6O2DYo+VnWI3sWbqTn5dvrg5cyZX+v85v59arXxlo
dCXUY0GwTo2879dHZHnidSh7afmTT4lq2k55NAICL4qCPRlB6uJqG5jbTQVIe8g7LRSQbGBskKOf
b8BMvrP6Qz/8H0Rxt0TH5f85gyF0CHNKiT8Ol04NtQhe9O89hynniItTB6O5Yblf+ysmLE4NBNiM
6SxOSRGSYyeESzZYvhiRKewJSBaTmZ6Z7PyfhEj+77qnfk7xg9oB58aDr6VHhn3yWvMTBxyRqiAk
qqI+L1Qk7MEBzE9+KI+l4qXwMRc51K3tsE+udw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o5YfGbeM/1z0RedW3D6OfyclCaA2vTggGu237RpCZerWjV695Uojlz9ps1iXCtE/aleCEUgSeAxS
QnWl/Ahwj7vtWh/43QPP6svC9/p1dQuFx9gwo1LTQhY/Vyg9cgzsT4L7i2d2gtGaCrhVOgqrNx9N
7JJixtBK2SAStMAXU2Q=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PO2aGz9jjKTIQH4LNUkNWkfllEuXf5NUTLtUhJ87ousCb5R6KFrvG8gZtQ4FRukHK3U2dxMST5x/
vDMd6ouqg8uNzcuEulW1aouvD25Gj7rbhPO3RziJ3+gRvELwFadUugTZsNTorBqARv21FA7ZiWwi
EGD3rr7DkYE2Nta2mB55e0jeqA57DPu/I6AfNkWFXtdQkIf5IiFw38lqNVOnUl4IN0rcVLiYfjlE
p0s5pW3g7SDIDhxwb51/AhQc+0b8to4lMUeQRsh4rzgv9uoPjBN72LTz4hfAoVykSM5OdBGXVymV
Kn3G31EWiguRta2Jb/US+lwgRty0Wrmyl3BlMA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74064)
`protect data_block
G2Oht6W+Knh7lcY1BZsZkGtjLsMiC4GQtDzeIbq/Ffa17+2CCRZjzXq1Im9m5d+yVhYljAR/s3ct
pO2OzS/A8O8AKIOYVlfcIUyxNCo6JgQKlwgJ5R4XcfVlG7NzXJhaggMPBr1NDi7u6bHyd13eac+w
qgrI5dAOKM0BLMoaeFbMUYBMUWZMuWCCXvxm3BDDU7WfzO8HKu6v/OePYgplamB/ZLQNLUiP8QG2
oqIaJ1uWPaIf8Pzn0cDnpFcg/gxNdYTboYUh1+yKLwCYoVjEa7zmggurdktlZaU1VXP50OtwgCi5
YmLpirAEJduByKa61zookZdc/8g6ccUBkqZgrQh+DawFhOmfhk9JcRq+xdJ7aVOVVUd8XcqJ/2To
r50XABLC78NUxZ6w2qq06bCXDTABdkeS0bJvg/tNKMTkP6k2n4aJXHhcsCplMtsy6pGHifx6Fmhc
MeKN55+qZ5HMWlBk5irGylRtgNkdHeCjgUbEp1I9Xjq+E0d3C9Lr7TZ9lIEYHgfEeXMd6pOLwzVL
WEAJnwImRaMuYLLfR9VGs2ANy3av1CDyeg+2XviKKh7/iTAZrXTEJV6jQCS/1AgCrYrMlYZYHUE0
BRXiM+Pw+zKy0Oo9AYyKNnQSVygDIm94Um7nRGh+omtQogpwMtYAhv7HjYODT2EKlejXNrzjgXha
6SzZJy2vgmkQN75T6CXog0tzpaVHCkctMyAoPM1YH+w6vEX+eJA5BH8i1qrKOVRugIB9ZhzKlIsa
nHLksJJlUj1PfXMety017d9HeHdO0Z50OFaf632INu3HWG71aZ9BhCesnbLTKA9xp4iDRdqYZZUV
HL4hJcTCX7uwZhde5Cej2JKndavff2uXN4ciHv44Xsq2UtONlopZGDiK2ssRei/KWkShgdk4uPQi
wxYRxinjDKy2snlnZCF7VdOyGk0EgctFcL+6wJ7SPR23hKPSINe9PUT0uicotnjDEn27KPlNFO6u
aPzCtuz3e5u+Xbvu/BxpP39x1nbwVEYTfrG8bXKVyc/KpY8KWk/P7BQeXTzhylupvz8d1EihKhMV
uKOGKSSIbZUquUKHU5MvgmynSu5+lplxdIwwlFv3fhvpUWVJ77p+pRXVIyFXDCdsg6hIZYAWy1Id
1fPcXTJSw7cKLKSDaByG0C3jVqtBZHVPJl0h4hOmYt1e2aeU7E5YpkmX3K8pf53jLYUIln6eML66
NLDVt5v3u9F2RdTBkmaBLw0dXHqkew9PbhYdH2UKTKF8bTde/j9qks0wkvQ0wN8SrIZ+1jDa8qBo
/fVxhUgmbMW0RFhjMhxByAYTkXRnM6WNcr/w6P3Y+xxlauuCH15Qwnh5I/rQPxgeaOC7X80Tk5EU
wIN2EfsPQ4C/2/wUYsZ7ZwXSIAzw6APjm5MNPLC3kjq6uv3inlQMwGRKh8TwzGVK37eECHoajsTw
1UvWWSF83smYkLpvA599WLLHrXdXdBvIfs3mRJ1kL2o7XUBSzRyqWErDaNOEgR0i/0ThUsU0LgD+
OY8m+P8rWiwBbv8M7jsDRmhi6eITGe9+MgQlA4Xfipj1nmeostiU8edumg2Wnw9SZPZddSQBNHFq
wdlVW6sgqBy2KL/08kKZv5kRp8p4VJrR0kJNKwsDAYSXbaSeSqiQJjAIpQdieQNupOoVGevpbtvo
/JE/L6xu9TUatud81va3st1ei36KdEnVpYP8oorREUtne0/Jb7L2/sDhOw+LwgptAqyr+96E8sTG
Zc65oVVGB+bzr5sYOWCvoL5V8SL/bOg2rRu7alw5eCifaZHXjKu0hK4qi5BCIoH1qItmSkTGWZlF
rDM+B8tUzFUTdKAdPHYT7hybtYZuFucB+uFQCZ1Fl6LyLNVtwbdSnIjmEboGP8SAeDLa+YT7Y8uJ
CF/gc5RbQ8CaORMmMrhgDvh9A6Vbdxn4RgAe/4+FsW/CgPCIkHsHkKDWkKfuBz+HKr45e7RFf2Gb
p+09NuuzgAaniOhTh+PZoFCcBRO7gahoSqbdcqWpw4L/bCfuBRCE1MjUiZ/olDWixTYBjnUEcInO
dfqu+VKKxP/0nRbTzrsqSA4W2BqEce9yZtxsIQgvvbFX5rgRZqPXOk0AvnEFIM0xiPtkpTgkSRCT
cZSIspZ6IBjL9HrIa7dhwQdUcnauJwUFVKWYrqg0AYm7wD9G9y120AjU3ZhjJDUMx6cr4d+reyx2
e7UcgnX87hjUL2wpBip2gq2PsK5A/rHDAqN40AugqQddzyui3thF9Upz5Zx6Dpt4Pkxb3Prn6VKi
Z7Xe/tQ8v2+deIKoEVOBufNcMhzrX3NWCsxmpABnXuq8KVAAwCqgM5CtdyrR3lipqwJ/BcMLK6+5
OfUCCKzp3BZ8q6yTCFoQlyBLEFIYIZ59jOqBQVXCjMVm6/F1My/OoRayZHHE0mig2ToBYmrO1bHK
xyRG9n7TDQurOs5xxddqFP1ZnWsN0L4TKor1+7a4+LeSc6rLMBD/TPoxaPs3jmfn2WsgU+m+o0Si
5UmdzW29Zhy9vsuhimX1AzX6qCnC5+Ai4yhBFYmBf9u9Vn3amdSCIiiqU/qxw4FV3eWxJyp7kl8O
05mE3acozDV3Gqy2LXuArWZPfAO9DNy9Z7ff2XKPRPpjsHo1j3kI0LkClSTvPmxRywtC6bV6Mldl
ycSrQlOhJrzA78QQHj0xH7DTfsYoDr0Km45OfL+/SQBCwe4MK6moxAqXSI/ZYnlZrJVzJFOHE9NB
hXA8kS8nhUOQVRLjjms+m7uxFc7C9mbcCGHW8M/jPBTCERhfIApTMUbQfiHLBfO8M/DUvVqfFx36
l6GeJUXxLf1kSK0lpT5aE40EhQHi4DzHdqyglavH5CkTnPOqNiemSP6iac9LFQWMCcxEwP25tiVc
cbYtgboAjolTSoZzuU0CkMjsOQRX9qOTy4y4QsLr0mWpl8Wzav+BNpH7r/pr+lzlJCtERE8EBMcT
mm1F/ehbZKhHrsqfHtICjBR864uRUqQZGMoWviApfURb11uQGGYjTUeffB67QvdFUNXuUJ5yyr7n
7Ur9d90BwQCVI9h7K2h/moor/oRhGIiOWMEnc1B0qjVLDhk8zAoYRHcrWqoHY/6fmp0KiGlQOOl8
SsK51e8UyOt7ZucEMJtzXqOmh7+g3YAHvfDi0xVzt4JPNe31CKFCk0Xmyeuq1cyEzPaZKsI/twXJ
Ezv4PzojU9Fe33/GwRl0G2vI8mdR2E+xbO0ICY5Hc8vn00Xm2kO83Mzm9jDOAC3RQ7im3Axr2N+z
UDLYb9LYtovpO3KI4Davph7YLSXPGmUaez9JFrjPr25pVKANgXU7fLwSQt69oqMToUXsBKT4E4e3
JBGOzCjSiFTyluJDNQKrtTULjgue13Z1IFAGZFSntvRy24af7pyaWNzGArUQaOtAKPApO9B6kAXY
ZA7gnQqdy3iPhUx3DcCE6UPVY0vlzud/G6vhVISRnc/4a2PI2u7JHgupjdmQ66bmVa8yKsYL7lZF
DSE9Bz/D4cBD1+pHLFWEtdj40Die8xAvHlD6dZhoOb/He50uUGxUEjZWV/OFJqJpQ62T2wREOe61
VyWx6j8hEql5Ce56j/muiHXBmYRgKoQtAhH4ndWCmbs4aei6cBR8gQDknXctI6wlCiB0J4HXq1ev
+wmvtqV6oEoqrl3+3bhIKZk+/kuhSNBFlgobFP4KFcaudYjIbCr23WAGxlVmz6846Z9DxUX159Wu
U5m4sM0CxrrTPHsGId6QYxRkhHFSQ97jbpxuGEjQYE6QXZXhLew563rpH3HifueP6I5qlQ4Vf+4R
z8Nh8gVxrxCRuLCQtUndAeBXra5NQZ9R8NA71OJLeS4xo55mKH5Olbk6MbBS1SK5UKJqccnzB99r
RwUtQGxLWmoQDnxB6tiJQ8qfxkVg2+G9XR0OYLcvvkJ5g7K0nuzg0+zbRWlEZHccbszK9w+qoMC7
TAT4RAZWZ0Hi2uNzmpc4omQOsziCyzt4NYvokO/FTOWr5wrE6jJsQoxw6FDXSUaYNOEUJDTYVXk8
jw8pOGPcwkQt2a/XCIMHyV/lkhqgWhDusm4eiRVaIfP90xoZWrv+wWTdDWTPTZUZEEgizqSPY/24
3GPc3luBg56P3CK4sgFMnTw+QGGQVQOFSpzUVMB1CF2sEdk6ZSLsiRfp8uX58akVuyZhOgYn2X8o
650oM5OtDIoJQBtj3grETWAMJitknbSrffKOd0GU2GeIUCndQ2+P0HtGpQPu0Sj81lKVoV3E7GBF
bmSfj4pUXc8ySqMOl+/J/FO0JlVaBbY3+K8jrAaEMBoZgEy41yhWa1nHi3ArT+qBpKGmVgdHaOG9
VmRYsnAnEf40HJbz5wZBCF0jWkW4l0NvmFr98RXw82PhmnDX7+3q8xKpVMorIBGC22NFdiFq9oRw
bL7h32oRpSD9uOYpX4dXBwewT4h1mTYVmx1fUHi/uB2MGlOV0mHoQGl6KLHXG1DRDqcip8B4iIvV
H9vaBC6hbwr0STVdKWKdmSo9XoC2sdWgudtlH4r8gjf3NxOMTrUc2CZ6sCWNudTa0D2Zd9Wvla8h
coLY7lg1jWuCQEWCGZfzGpPvi0hC01rQjMfWUy8qirUMfTCCsUyGdGmbzuxe4HqfSDGnp1IMclVS
dagfCO1zZ9jbaRwch1Ez3XRkxZWitbnvl0ecuDhNxN0qgFVfLUbMax+lq3pmFYzw5CpxUhsDLgGW
xPsAPoZAFiw76gPUXHvtHU8qmXOAChM4MLrbhA9sqVCvkxraEzijyGZTQEfTUdYIN2TUqJEhc67i
MqysAj1AO5O+fZ6RrwP2BHZGS1gyNIP62V1VuyMCQzY8RvOnNOs6/OnROXF74usF4qokK7w0/nWs
ZCqFE86EeMGB4P3Ryg8shvsSeKLxcRUaWcuhqa0CQiUj9NNDAqrI3hM16xvjyuOZPEt3WrkomVk5
KiHiK9iwVrT77s+c+IjpGRazazXG+72HmSDfV85IJhK0DuqDcIHMtUVZjdpHO8dJiqPMAFahlXOT
HS/lL/Cox0Rb0G8zot/diB96gppC8klx756Z/wo7VtYfCE73L56pm4fjaTBpnWx5M6IXcw/Q3BYg
UTjDZG9HonNcyk2iauFw5gVPrZQDobUxe46cr5uh7v348oTDn+Qg8hpXBhsBAKMnDSK5xZGtkepY
wlxaTNiVxygWqCtkunohX33PAYzHW47uDNtxoWlwCWQKaac+5ho1GtOf4MfA60KTUVxyArDoDqF4
p07/QL1IQgD5BAVOY3mlSr/mGlnEljQbvElybangM2OExI2FOfFU6RqlfhWpcCaTwN5Dzt3JTvXH
owaEpB/U5K5Nv01eEhg7YZZ4Fc1sNEhAFEeM6w892jtb/8ULwc6Z1PzzRqYGbc5tBaiQTI/94mC0
11NSGfQ5zGNoS/5iioEKo0mPM93MqSQ/9t5QIzgjcAinZz9A51+S/F37maGwJ22Lp+8XMXiMBhF+
HKJDplmGI8+QdpxY+XNlthV3fX0+FSyAb8tF5J6AtrrCUpHdd4H0kJy0Bd5nVrNgi4qHyRUzOhRO
rL5zx3+XVk6+wsMVy4vvNPPKmy99LZUejbMjWtfyVEQ6OnrYwhRvFgrcwMhiO1lSaYQxjSN38Ypz
Z+2z+3nACWy412CEqXL4YKIF1u3maOYAQkb21a+i+fPEKUdznuqjWA3/pBpS53nN/I8wFDa9oeA9
M+hoQxIMiKxJX7mMYdfhHuPyFeILDjYwpk5OBcjLZ6ca1q8h3aJxCMMuIPrkkBtxv2acSjM5SipD
qFxuMF0ev6+2iPJA4auHIYxab3VPA335FHkl66hCVGHIioJvukUe5hT9lxz3wLO2G1O6zS4+rh5L
/+GY/onGsx3glhnMxlUFbcz4Be7yOQZ0kY7aTJYXbO/5XvmPYK574ogcEX8ngseKKxY9U+YCjXT4
MDSxX4iQGGYw00ANb8Y1wpvwJ+gsvjkvFjM8rl5JIZKwt6S10iZsrHM47MdjCMuhmu5EmBt+R5Rf
JSQ1jZxZOuZxqog0tvot9+57knB/jt2Q5NVyQ7nTGz6Mgw6QWDLj5QBq9PJgyVz8/8kz6K8CcWxO
aWrp7qz44/LkJhDJU0vMSnLgMGzXMXGxIXr2/YsHxso04CbL/KgsukmT/uZSCght2J95GJ8WY33S
XDIEr5XjeYnkHlp9YPQ+YR281KsPxGAGsp1i0t08U0ZXeNqkryyzNQ4OzqbEHNCujZFR2Plc5kpG
3HTmiYH0f5fNA5YhbtNFaAZ2TIP4sE8QBfRDefvw5YGNQMQhsBprYRIeBmsvAHlUtKeCRRrIXVn6
I/neqmZuya4BUW3XbAj6u+lPVW7XWvJi3ncMjhI17fcRT+RJIXdhdTjyuQuabUUffFO880cp9/Hp
8SyhLqrHTXdM4jf05Jkss4qkK0lVf+2vBSIMB5z5yvvamaJJOqaWHDgCgZwL2cEzQjpE3IuJ9IZj
qQM5kc5msBYjT10TtscxBm9MAZ4aWLBL4lfgrOEGfbeFYQyPoeJFiRbCO5MK12/cxxCcy5qqSWyL
sE0WKwX/YJ2E59A4/kgSYuYytC/RmqQhhE8+VoPnR4T9vrJ7hos/U5VajfoppQVVmR6aiJkq7VLA
QpHjB4O0MoLznf2tnDqLBkWlXbeGcaLrT5n5Gklvt7hdO0qli63rN2x2VPaE8Gu1TR2ZVmsYnHsK
qf1HNIJfLtd8wcFtHMuWe0on0msKKRSGxeqYv8W2QF82eRjGWaarNW926sEh1kFtjKbXuXXddpFs
lSUw/JzsI+PS58LwFedteF+umDT14rV5/WqCfkwLd9zVV2F9X7+z97Y5vYx6d5xbHVFbnR5iulDb
TWwA4pnibhBNjMAO4XwNXSAhPoNCDJypgzfGcsxztKRn5aqt3mm9V8QtuyfTZxo++LZFJwALuTEX
AgowDYHrqBbD5tXcttiz5U9OVVWMfhdkvzGdDUFR7TpzZkHM/l17rOymeibCwqZ6aSq6qg/WCQJ6
2O4KJTEMQBbXhHf/1ghRkVIrT0Cx5KzayG9hUALz2QJ6g7z3PVTS9jdyYHBj9WD8wXpvBn0kXe3y
e4v0bhLftDY89u37YXQI3JzyGUrO+cyR5x6Cm+71B6I8sGkw+wlyVciFMuVnnCDPEhsla8Ej7iFF
ZAqlNB92EtjGKiUyDlNEyK+ZrQs4Nd3PY597nB+o8+DbVeWRAJlbftW41D9ThNpNMwD46O920+Bx
JS7ssGdWVf4C/CWbjqCM0cuDjwEIMS7aDzvniRqOj/ZgJCvV6EOIm6nep4SdBfoReTMT0ZxSh8Ym
litFXnmXVogRjoEFLqeAfwBZXvJp62Fq+/J+PlV/zcto8bs+vvW+FO9JKHJYscA5v+VvLENwWt1+
RDNQhfLzBRKRAiZx+ThOTdtR6dymx1mhO+CU5mW5kLSUaE0V3Gb358cwwiiLpvbXZteOQfEANEbX
eSduZgKcFzTGgAhtDU/eQQAAdBgDRznuAHDcUqeCrTMCl+d08SgtojS51Kz5YfY/lJdKZ+J9sQs9
zsiH7vNFeg1HBeilhMAcB3WQt2QWan0Dn58R9dddObAV9G8dRlFqYX1OxsbVi/VU9LURJM9OUtn2
QY7shn4dLT/oVijOx3kGVtQxD9mcz6sS1DDvwKZV+uqc2RuMlEtllU+wO4MPSlp27JlrdzjRyhT5
+j5NCkx2q8FreLYdh0Y+cnnYDxv/OCdfLPmkYjQf6aJQUuL7r7SYDi1vtcczlHrrfhUQpna6ASMR
e3PYa3q2krc9eDJ3HLd6gdCc3DaTi4oHWA0jnbQ7TyprQlxa4ETs33CgrHLcX2Z7xxLZK784hKVM
6qOyTKNjz6gY4jltuh7a85fam6EZynCiNL6P7MaqY3QFRHU2UVMvu+y2LN7kyerzjGpf7xqe5qCP
trPpJIF8GfVbwbk/F3IizREU4o7zkFwn8DBeJEIJHtZASzaLAwEDmSvYbkegugOz/MGPAyQpNP4C
NHotxs37rC0sp+KfOrpzAFPkX72RtgjOxPpSMZJotzAAhwnBSOM19LtQRa1bpYSYSrWU5WQKBHBN
9s8wabctjf+l1z+Kp7KW85/UNSrKqvUXRbI3CuGT1h+eNJJRjCfQplddofccmhYfEuP9bX72YAM2
Ut45lXAYaNqsXztFQsobS74INSGNASE3FuXehLHCQXhy3Qvc8fYvV78oafpSuUf+RGpo0gCWHjyS
OxCuEl1Tpb5jFP25FvWi9T+lFuJRcqQsOalyMbH7ZBreAv7aWU6wTO1plGOiw8FVv3n2+s44BKRv
pwannFhgdO/EKl95xM1okLy6Zf7wabviGRCTjbNSyL6JyTZ0VTrLpoIENKLi8mYWyorvCgYpZl+r
67IgUyJ77y/L3JzAiH8a6tKZMbA7m1vl0dXMw/ohJoKTeWQXxEwtr1nmHVUHm37ySUZZiw0rVbpP
NCwA9524hE4ToWNLI5g5s2+zuxHMO13b/8PwF1z8TDRx2jQu9ZReubWQNKBHJNkNuolvBXeJ9b/X
gsmcZWBWqQCvhvc3i++Fyk+0+9llGCglZ+m+y1Z+VigmMv62YlQpyl2jhfY3PS/+77awhIAXgs2F
E5k46rkb47Txvm2uY758jU2GdnwLoi/MGa407hgy06rY1Dmn98sd7RDsy8kzLzWrv2xHPplQ9pSm
e7tS+zC8Sg6oDuLHTr1zkY1usLpGmdNtGica34ee4gWoOnP1ueUzapvcK42sXmQWCMtntJkraSo7
yfmH6YGgJ05pKsq9P5of5Isk6meB0n3dJHNYJrno5nYHSRWphCWmdTjbGgATDqkn9DNdna3OjyBA
GBXyiFW1iBrj5vSuDotjnZnNBHaP/kSi5M6RTZXyYqjioodwoiDoUPYv/DdblOt08jW/sArKPG7T
i9Hz9BznLmRbbk89oaCB/OPFNARLxRfi43Qt+533qBsAhxVwkfkwjqdDrrthHQOqfiJo0gMeUunq
9ddmg6mT/P6/+wNa0LQ+s5Ah5LZJJdFzGpaqzqO8xbnEDvyiXdet+bytmE1y62zu2nmeTNmU7TWw
3fiYksu9SR0K/f2V6XEnMTCO1snXPfyeJgXzQFpK6MS0jo/8/q20zAAR1KuFRM5XQq78MgiLggHI
9dRQoammG7i0G6YWzsDgZF6pmQ3Fb02akA5u/9YzBkSjm1UB6h6OHy0VfHMmmyDBJOiT1LDqIhCC
3eeSm44JLZQt8COS0xNZjbLl32b9nMmD/VtT9R6yv7hQbl7CXc4Ii9n5Q+kixcgNYI2eWuVZzqKO
MTCZpijs56TS6bGYfALeDsGsXnhqvvgXwtyrH7cBZOlaeaz5LqCT/b3wfaWLUJfG0CEWxCO3FSDZ
PcwK7a454Lg8dgCpyuV3hmX0hkk13JITxPQuy9xl8rNFbnM6V0vPkL67J48LinfQiIDmwHVlJabl
h8QzXswTBU+TyoKBNLQQcNjNF0gwSCEMziu/9OVtxTjlbs7ThKpAsZ2t1+rAsIKoletSKiFIr45I
f5ItW5M0g8NJT9qBGCxhmhfZlpbu5YIVTgne5hI47IjBPVqaOSazSGE+uEIPdYdWtDqLcLllqgXl
xsR4DHpkgjrF6sgveP7/sXdwAu9ixLCIJft/Z6WzxlcperPiSkAQGBhhliVWY1qJuv5POUXcIxZB
VxFAmY6fbEXMOf6qopF5aAGNUaasL8KOvy29brbLVBsCeRDtZQyXkgo05KZ8c2N7h1fg3f+8i02+
sBBsUE+E/LJ4wqmy5tj4umbhUrWhOzMF13K13n8dyoNe9SH1+ZOH+FQblJpkhwneVX8/pbW26zfx
o/K6/1iAU8mBXT46lsJLc/oztXsYDmAu5r1fFqMLvwjGiTas8b5jbqUOz/s2x31gUV7F0meBP5vR
dTeB8QYHEFqUX2KfWz5G6GpwWprk01QZ45CsYc9bkPlALo0kZKu0X42SX9RZfIVdQogVXQhvplpO
7f/RuJ4eg7EjkXNUd+WnZhVrianUQ4G+Tg6kYG3pmsj/Q29+oNNhIA6AwXd/90cBGcJHTtpunmUU
+l6VVNnSmq0yutj5qHAMOQ+Af6rP9eoi9LFUAMkkQtsXxzhghcxyTRaS38lNKLRhSjTID19/0H6C
NQICePQ8DAnBVksWCMsvEGtHqXBkcl6i/fzIJtNNxdYR2TCMDiPrAmE/48kbYmru1BZPKD6cO9C5
7sIh+uyXoKAzdphnSjRmX295pCj3L4sIJIN+xzMEYrBb+m+uBueIEZbh7aggRhViQq0Y2fKyON9F
pBvto5jVwwn6C1LhWkAyXeWOkUxDddIm5c2vSK4sthbD0eFAtWroBER4DDqylKYUQu9aWyGkri9d
RJymcTDBEuJzIf/TCcg2fMCpURO/LYmESAx0zD8fQyXqm+s4Z2SCP4G/H5Uv40iA4F9oWkJlWUvG
VDn+t+zYmqnXVTR4HbBqpZhLcW1jhkYGKxh8D2kbTtip6zzlSfY/jncSAfX4PVUzzNZUHX1g0vPz
Hqn4M/cvdx+mYLxFrbBmw8f7KOToxnECJ/anwpi5parGLvTilCZ2RAfv/mglhQK45vyhFjgWwyA3
hilTnDz07uOi253joXVv1oyTOGiLiHY4LgW/1LoDUOGTseJEeqePm7LVd/C69BDdKS/kbebQe4zX
ozOGJXTjHtj0b6J4a7nn7ELlGjKlA1wEmafUYwqUc2ZqRAR9hVOC1ooVEFh6ZsIz56CexLCwV1wi
6AM4c+G42CsUv1WLQLdlMVZ+7AprG7xD9gmf4rgQtc4OO3TcUYmWUecjdEUjunECLw7ItslSXjLX
6iRb8W8JAJtKMxRe+7Q22Vwk5r/p8LFnBkIYEWQA+EbSC09FAIhPVtyRQS2Govd3CEYlJCnwBmL8
QJshQioAbVV74VVOite/bZXNMzHPngDFBjPqz1eT1tPhZCi/VsosfwQryyvStMffh4Wkk+b4Uvmq
L1HILk1euQkK//JRpDu9QX9QeSEtXvwd+gxTzHStELhvTPMoeN3taaVn8dMhsIDUoTvTKMrXsqos
FO7x6LomX3HWtJXhh+XFT26GtffsX4ASSPr3cg0M5g1nwvH3SJjdxfVkEHkOSSKp7DiriyNjMnen
EZ0d9EpLTA5c/d4FkW4COyP9rdTw0GNwg44+rZJBUCFXv5smerKyI2kmAwmluf9dp+ErNY3WrF88
OM7V5X+wNWbVUjQhhqCSnn+HHqtd2IijxZMKpwjsOXGuIZBL/qj6XiJXr5bqagDN66qioMXIffzB
ZNyU+aNp+UdXHzVe7oOLEljmIqMd11RphHq+o1gOhjzAYRP//aWed3g1PDPcd/2xSumFjIbDnZqB
ysEIaKfhErmRFpgaB5LCj3Gce29VmQdV/oy91/5hCbw2lDz1g0E9usAOp351j7sBeWq6aiREc4S2
c38qJHqp+zCp/SR1tiZVYT/ZKDvrIR22+t0Vo/Qf6kJdtLB02eJWsB4y2GOiqSp3ABNCDMvqQF0d
BoX+1A9rq9hlfDyx9FLFNLA0vwpRyfPaR/TKy8BdB223gacJ31YaPRrUjlvc/UfVFBDnuXmi3wfF
0VyCNZ6XA7rsyftMgT/EQTC7b0BlgFOkbHGoIAh+V6nw8zKha87hnhh2VDipLZSuW/mifGuo+SZv
nOJTss/C/lFxmQnDV4+Oe4G8KgoO0TnEBKrfIQiuboa7sSOTtGSgprzc/FQMPZXoM2hPogUkO7Ol
MjgQkGCRTPRCvA7DtkPS0UmpPKaFfUlMSg87kU0RCRMwu0qQoORXb/WsK1rxWXsn1N+PVXQt+aAN
V+pdHEaeqyXB89SaSq45vZk4JoISR6YUBTq2Zk/yawiM+kMypxHTzlwjfyTkQMkQF0VlrxvkXhGe
7GFRE8fkb4Lisd5ysP/PufbFi76yzRyYGbp/Q+H+CrBgvZPAGjeqFgSnCuA6tVCiiNn2PEIqDJfu
RTLehdNfS27x6ctv+dOuaUXl1HpkazLVcyMMYFYonIvZFW+tfpS3sOyrSApw1RuBzwr0wQpRpAx+
1N/4lQIFiVVfE5ahgJ3n2e3S5n1Sb1DweUXwhRj9vuHmybDCGys0A4Fg2NZUu92bJ1Z4bIT+Ffkl
ykmRE2nRnBIpxdMZAM2iRbWl9hesmhxTa9NuODPDrpek27NJQ7Ub3UZUQt1QCFrmjyXAFkZFSVR4
DUWwUnZGs3pTwzBrwB9TF+LzfiWyzoE35nkJ8Gbq6QbWKN+WeBqE3fieQY+A7rXBSqRyf3IwJWG3
jmJ/QPkF6i6WQ8ZU4LWN6dbblVBm9woL8RmbFjbG/opxRYQFA5o45WUom2aki8AtT6nDsDZVbBcw
mu/yk/Qf+nOhHAzX0F9FjfJZk8cBwKjPNoc5J/WXS6thl1PiTeaAf2B1CR2RnOKeXT6Zl8M8X45i
qz8+nzi3h+EKCCuFdhc6mZ2+qCYzrksf7HwxQP72FcNbt3YZHiL7nTkjYQh44V5U8YfThX9roIoJ
7CMsfodYsC4XnTCw6qc+TVreW4jDzky3hZ/xx0owVXNWiyr2u/UrXv2OPPNCAqh46W/3Np6AW3De
DI94WMVs36T7AfvOlWCyUvUTMrqB1HEooosyS+RiBHmrAi1RAz9HQtqKUhgHhX0oNT1FtQ+mIaDn
PcO6YuIOHUqOsc+ev2bhYFzIHKV5BTM+5z3zu2Q37ELK1lW6MY4v5/+4cCaeGFUI9HgekGNFDcC7
Hbj3TKbqCGY6/WhNzm3Ru7XpAWnVTUxlQ+BkTvle56reilfsvhI5WYaR2M5A8E1Y41zZ6gXVacPF
senWq7iEoqdnL81fC9+3JuwEqLS2c6v1j2TG4Gc5ZyFf93uRhliYIHU3xAWU758Rc/fFGsx8Ah/H
FNw3MPCcs3JcBruvOcNVjMOA37HZx08WE31RKs08nGslcwY3R9Y4kDXoFqRoKG3MrTWgh2QqLgv/
WvYuKxOSeTlI1ixYGUbMurtxnD9m+Tp3k0xmu0XIeJ44hcv6iPkMFbprYL3nUrhom4zgf4CEbPHT
AvM0bb4u9djGlVhZk125c0n9DpQjg6e/sf4NhgrSZYPSds2597TKpbo9Gn/jkvDln1WGpOeuGakW
ZfNZ+g1bk9p7Vu8tJUET9dywPBMpiu0ahpGiXug+UGO7hQRWNR+e8DljtB17KKxHp4aSo/nIQalr
afh+g2/dDqc45dHoqYPXUHldrARgqTNbfFwVNMd2BKuxtuEGsP5Tcd+zzV/zyhaPZ3OmCt1upaD+
1yxRNQL/86dDbBxPamvLDBS9I2h5uVGqNGDaLl4p7dMA4/2C5S5ipUMJ2BXBdfbWl78VvWk/K2TC
9m+ZWBSLt3ZO5lGqmo9T9zzPIukxOhZc/VSnKfsvx2H5DWC2j/461lazVW6XRbnSzaqFPSYOrS5I
BHvVneGJfcyrC8K1HF5hqW8KWU/uB/P4pGzsqELD8GkoRrnRuj0sWD/tOcaoAW9R//tXjVSGLBZL
Kr9Y+VETLkpr/uBgFyVazAf0437JFIgb1xP66OnVskKNZSEJg3zNiEKXTDHccNwTr6XSFFb0vOH3
bZE9V8mtmEZE6ERDtaJRtjKII0QZOK/9u62wlLvEriunfBi4F8hQG7S9bStmY0SD1eM6YBEP2PpU
iRViQmCkv4pMXLFKtq+6sXoxLX+YgxXjHuBXRIg5a20FzVKTVGZTlRVOLWm2U7hkSI31dmWHmuZB
/FZQtWjXL2LhriIcyP7jrG2CCEwqXzDRyGUN8UuzcGphuuIwSJqhNLw5buC24V31SqkmZbmW6U7F
cttbodh0rYuE14KuwjaoCQ5JzwVXOhdtEOs2v7GcMZeKROw6hyOiFh5APo2HAeLaYLmMj87MQYVF
UF3lIzyTRCVZE0Mza0ClkRw2UdgPcnq7yaZfS5dLGKeYs+C4EBCb7q9xQigYpngHvZa8rNe7etBx
RDX353VHxAkyMnz2HJ41vzoEPW+6Q/CLWUKBDLpeKSI7W13udMX0W2V6CWFohaGnwfFbtx3tesJR
1FvIr4SymB75AcpeBQ9vsiw3Jn1V8O6/sId9rVQwu0gs8Oe1k3cf/HttPjMNv28HKHphhrxmxtxl
xCZaGzHJFWe4oFtXGETbxeuo147xXuwldM2QyN1Yppoy7Jr+ayKhqsoHaMJm7ynQ3ERSwdyhz+h4
b+fWHTUvASm2CvQm5rL9OksiuW2QNi+DqJtdOT54ve6nAQywQX5IoIO8rPv1gPZE6kYeVAdjQ1Oe
Sb0/axTga/Lf/fsqsYMy0i9o7QMWCHcon5voVmLlKhMJXV6NLoIGREddSqdot6X3Ny7MdwHmmfyw
ycVUyeRrcxLUE7H0Isx9TWezJGfcHIIyGlwMl6XJ42ThIbY3hznEcI4IQkh5TNdZTk8s3p6iLXjL
fwhSQHdaBN72WMM8cPmeZtVIIkDvEDxuwBXjFWu90i5rLb+sNgq5wdvL2ocMLvbryW2/GW9foBjs
AHCd/SPrK0viHBcoOsDa0pBwXNkm9mllk7WjoAewDjgeRFzM9e6ZvkjxepsDas6bwWS+BZvz6clw
CN7SNdbnVIGaux93B185Ms0IAI2Qi6NyXsFq//QCiq5XM3bI38NXqn0yda/DJvli4hyQaliQCJML
wh2xborhH6M44Ok63FDy+6HoFFPMoY4FY819u4JOYTOmiyYuzTih4szguZmD4kOvauh8z5eLfNQr
qpBosCoCaZo7PGMCnbgxbAIdcY6NyUHxjHHQExWw6NT6fs96uzRA+dC/c1lJ53BkgQanKx4lU34L
nScdpRauE0w3pQ04g4CwOHtEq+bBfzqx2A4uVZmLvrsUuZ58Pk3mdIbkkB+WUdPCsxpDYmTkU/px
VS+bzO5Otxwr0ikYO7+49LQloK+kY3NGQ7WdmidEZh7X6HeCtRLYM1sbygAPVpWcjnw8q7E0xUkJ
n78wpyOdKkc+j+o3G/Rj66+oyoA/1qoSVtFpQptQs0pDR7QS18+ZOg/loQMzqii5/58Lwky5sYb5
H0xL5eS++oczJX6pj2V0Zw3w6dhaxzMEfE/Y8da95flWf1VpNg2WCtmLCCSGnDxpMemoVi5kzOHs
Pz3IB3u9Of6QkrNA62J57HwGp8KBlMBTxCEYOHf3dVz1L1lSYb0Ilh7BO9eVv2lfGYjpZvJfarYd
+w9LgkohX7JsCFRGNcnxwUGLEsY9Hm6Y3F0KBKo/UCfvouwOCfR0fZCM+c4Bx1jdfA0zvbSDayYA
jpNpheFdkUta+epvtwCNvrY0RUykiA+42hjVeAtDDgCKNkuXguNeXru5HmJYmMuc15ucf42F3uF6
tB+hz2zvn29/RK6Cdov1LVboXYbyGzGAHvoZWfgAKcl9HEfRzg5K5/YEW2hG3aIhOzMRAZZqg/iM
YmkJgmVNIT3luOWWEv/FTq0TxF2UH8eaRcwLL09QqhcIorK4xd5ACfyDwX8zpExkKUczRIT/gUOD
BajAD0GM2t6J8/9jqLY+wKnBELTilFzqm/uzmOoLoy3Z4TFLy+kix557Ba1q3iy5O0f7IZA/GPUr
xTvnQxpWbervwkelJZrG6gYYeICzm9O6+gc0FuNanbqyGrXZ7OsneGVhnepUUbHgg4xlz/D84KOa
Eujpo7eyLlG9cz6h40Y946hNeOM1gYIHNC13cVn9BPnwZ0dv6K2EqEj/LKrr/it190iE4S3cBtOF
0RD1IQnGEcnl0scB/rAvD/fTTP97A8e1qGJLiBGZ/JvA2YFqo+Q5b0DVm9IIRCWZ8aTd8uSMap5I
tD5cSHf7fWQv/AljVOhoCQZdgO8aS8myxYtF3lwO0jwa9K3/HRA2FvrepflEoaWGgLIgrY5Y2bt+
FLCYtu4XOozgNGsrjAEVVNIGO8i+IEqdeniEXzTlFvKlVa3JKlaXLwP47Z9g0WFtfTh65BKI1VNk
iu6TTZipu3IEeXC3Q5ITxyVMqzmGi01T+g4/lNKwgN3rSH24Mrgtv4LDYlY1KRKapP8e1clPeFi4
1UDv4lTcWrxp78ZuVMhusYVyCqdTb7CPCHb7dCkLwC/nLky6rFlV0bnDLssZvy18fc7wkBfCI/Fh
8aVxZ3C9r1EAZyMzBoHngWuJ6Fq0h8A1LFWE7Tqt/sr666hjffmyd1pnwZDfmbwBIcNRi9GS+Fq4
/6q6ufElUGfXJ56FsoL9v4qhrD2tyiczVnljFmWUl6v4cy1nOB74acOeqcgxSO40FBGOiTG3dbCV
G+Vkt3N6gUJ5nNRA1NczsAB+XqliKrQ91z8+kY55qyYobNORoKjcBRz/aI9/5ATnraBfRHX+fuOD
Molhpza+ngf23XMealBnWOKMoOEY3m6Wt8ZWrZ22eGOd5SEDAiUS17STRcETLZWGSde7GhiQQNsL
1/kF27qxLAi+WvAaqIJS0O/QleCHR4j1yukqfMFQYBIe4Coij4x8Qyh4mj4gNUoT0dfoD8gLoD1I
ptlLS/59s9FuBuW3rI8ooHFqn/GvPeVVmvHdPDfIZtLxeKBcuIkCyAKpXAh7uW620lNufyM1O4vh
KXb8p1jnsm1Xvmk4IbFDxj98nZtXFBmY1tBNdFTFweuqkK5b/Lg2mvsgKhX5HjQHUfQRe68tTJPk
urJDVcNoJ6DUJ9iRlBvBE416BAPsnV6qGEnYcYbdyhF2f3Pf5jwutgRYvm6iT2J1uX1Lx6yK/PMj
mhdPu2xLTrih91WyqrMJbN48HKQsGOwmO6mcBP/Ew7ETMdEhc4hdmBhGLDYawA7Gd/Blf/1Dp83h
jWLOPUhvpyGfoxsig2NVkB08n1n39UeAN6rsNV/3U6rpsFOWPjOUGfAeFL03A2i+GVp/Vw5oku20
RgNnEzNGkhMEI/WKH2/iJXXhtSatyl15fciXDE/n6WYyLcYoQ5qqC06BInz+4e7UgYUQMJD1Hrr/
ajIXPu9BVl+RhVORYofXEltLOAjr0THXRi+18xcMBCqcygaJa0h7z0nW5iQjJMG3fcg++Mnm2Yau
hPGNp8RvCQ28zt9IjPQ9Mvz6Yu8b+ch2hJb7bqas9dziNm2bpkxCYXcxxh5vSSOoLFw9E1b/dqr5
CzBilzER7vlbeRy03UIG++7ILOuE4EMOw10Lkkb2uKOlr2vnPxSWB62lF3CcYzIQoMRb4AhZ+pXL
PZPmDEWtiTnjHfp7VscE6kmYoD1nr34ATtBYA0t2VXBqD01HZEPqK7iEksDWR/pptZN1QhS5ukAZ
nsDEk+NMhnQDnEIaygIgZR1TMyo03WtwebAr0sdFqXAlctDNcQGjvpYQScSG0GbF6tDmvj4FWLyR
dukl9Bu4DUdK+PEbStExqSaxsapcp1z+vub3XDDJoumXA+SuMs6fjuq6UZkDJCWMXrk/CBmvQ1+Z
9Oc4X1o13CrzPtJCeUiHn7ik/sJJk784grH0dZrNdlq0osBjJ0DYLjB/iyHu8T42gFBBQ6Og/CXO
hZYYIu/tTbdWLCViwAw3pY9lnX/scqOtv8CzN5RXWx1rhX2huW3RT1FJTwPQAzzkyxm8bX4O2cs2
dUeSZISzHcvJKSrHNZIsLP7WkmEqT2XsVP36UBW1RnWvvVjowDQk9uk3JkDtRkD2soiOhI09qSJm
LB0sOn75zBEs0/cxd2NUemTkRdDMyNJKCbn9Yv4xgUqQBA+JTC3n1HXoDu95zUE7wtvWVTDJu2/7
v0Yq83v1uu+TNewIyl7NMoTFC3b/xFxF50fTAO8TLl7zgtbPcVFAT7HWoOn0hFnHoNKPHREklO91
8dupH0lgoHDxEIGZJ/ZPhSZ/A4rTVCrXFZyqofQAw5GBTGKqekv7N8A8UgY9JA2FZXiaIKQO1Wkp
nPgwCdZzszMU9hx1fZAnKpnip7AwZVEmq97TTjnhlnbMDMeksMm034E7npp6osI+dpJBujP9uO//
gKTO6WIU1881cxHRDWI0Jv52J/EjHMZmarSl4klEYieepwVWbg2DB0unLFvAVelIoW46ceh2jgjO
TzUbE+gZLEKp0bXBqojeE1RpDWDUhdT1TEidVvIm2wtRJqRpK8YiMVozCe1zAg/Iwn5FzSVcqJEJ
ZzCe9fmQiulzWsbc4Ml4U9MXVDx2wO3Z28lZDUeyWe6zdGF19OpNOqzGeCX+7jVK0ZB4SEOeaLqn
UGE1VFVlnL6M7sN+0zrbKbcNnZ9MGx4peqPgNgZ/28Xc9o6EQ6n385KoAhXzSCK1dMY95Xi5s4Q8
fYyVEbms0NuS+14K2tmapndc+1DF3AnnkB1oANj/vz6MFUP0rcv5jm6RzQVO4ZutBA6se/EQMLZe
qSfEzdxi/u1OyYBCiEvMVk4QY7EH684KenmKzSiW9vBQoMYjzmJsSoHF77awE4py8ATaMfgqPLk+
15IEn8p/Lo2ZH+cudhGU21mMdrVz5QDeX67Qta2UsUGbOkpdWajAAE/iQnTwKZ66Kn7SrWItQzvx
JmKeg8sqULhOyYjjDSpEO5C8XbxaTK21vh88qYAzr7uSzmV7ODrs+VZDpCjtqZ64fFWRDAKwD4z6
NoOdIhMk7Vi3rz4goL4Tm9V1NLANJtpmYuVGqFVM9PBqq6yXj/uTiInfGEZdxtSiV7TWNn9550OQ
w3kbeFAbgC9wvzCb5rhXRIbDwVJXD3SgjMwHpn0QmBnbOgMZq6u9KBvhz6+S3a5pTwP+m0VeKhdO
rZeRC7EkGVeJVjge4mSF0webZGOkjzaectsFr3K8OQwHXT1fvUzHRRkdvRiW7ZPXH8PYq52zAZep
UINjuX9u0jIZBznsVXP1N7ldRiV8a3lhYWCXCsxpQjM8nyCtTUOOjB32awpViwQl8TP6nuF0FaWq
J33y7uHJN5vVkSRfsRTXyVNdSQvUm/aZzfMkiP2N/Ds7+plhwfsV3WtOLKpjwS2ZfoMmx7OZD7uv
f8FwK18bF4m1BaUTZzHv6URcPm1bPcXx9DdFbuUXkGzVUjtewf7uREb1p1wlRd/MS1V1uHANB1M3
gcNLCFpammcHRjWaO+w+3PrV1Vc/tj5lba9HAH7oOpxYgNHfhRqh+d2L4hzMg4TQmg2zVglP5H3Z
ZEXSHT07eeWDOgcZT8013turr1ODA6iHPp2I66/L7wZ10UNxV2YmMcYPtUPCs3A1wyrBe6u6IwZY
5PTPm9HsmAAJO/YMd7vdzPyvHjZS0ER3t47uRUpZKQ2WJu5dP3G1sMmvw+EtXNUN8Rw8hqCT4rXT
aB1LgQX+8mhMV4tGJjCPBIyrQqiFLGzAKBRVAUerxO/pRdugEM3JCY7xVDZ+DtImodcwrq6ThPqQ
q2MVk+teWwSb4KA7USB8Q0sFjcovSJKWlP84uFSZ0hL/281/UxpkXw8Wheou9h8ctwMkVqlaH3c1
BnWXj94b0pcyX7+Q9lc42Q0UaYtfUI+R+sPqAoosdz49080Byhi3Wf4sJO9H3RojwZP3JPBAKOyD
e3ZBPnqhZX8jVdU43RJbrcf1SCLDAlKBr4gjKiNsI6QurOXi+gptf1BoajKj6uOB98KWeRZ/jnqh
jlFRJhdBlTAIpByG4ZFXn4W2OmAd8D5/MxnvN2GGLtLQiP9OV8Mhjz0hsJqvmf8FHHVFyNW0xzr4
dOXeYHpMVZn/8QxRpj1xpnoEZ7/VxwqOZ5THwKvladTwHsSmFiXs4PfHOg+xKA1XlTucJNf48/xR
WSd/N82FU25ZdqYesbioFNUQAR6rFy4doNQ4Pxk1Hk7nDdfNofTvjN8aCUWx1cxA2nPr2vzY1pHV
JH3eoGpvW43duEmYku8zRULL0rX7iVZJpbmW5pbp87Bl3Gh5pc3R4fslWYczkdTSkSMKaUiu7CT2
WnzDC5KJprtBPzZyed6BP4zpJfKMN+VGKCWdBOK+pVALxSpArqRQmSfcqTKJKM/rlaLXcsT5PjEW
4hOdOWdF7q+Bc4exgUR8CGe+m/p6uy4A60x0a+1tZ++qZyOpxo9omT8BP5bPfwZqAXC2Mbq0b4ou
3dmDxSCFnDi92NIuPpkXahL9yYy0xCbeyHDfe6MPsSO0uui+5Ou7gyXrmratOLoG/TisB3RnO/sw
kgGOUfzgzf6NREsS0arUO8Nvlp0AzkpTeWxpP41eMadYguGz49uZGtKz315Skx9bJqGY5BxiMCcx
T0DkK2WuOpj6xnww8ibil5eX/vf288mDXgjQmeDJ3rJhclU+fXOQPe8ddfRme2C7LFfkICx+ZT5x
3EqdVog3OsZjln73UbSYYoNFOnowDEEI5Fs5eJSmVsEIeZXCy7nLf4jflyXM+YfQpoL3WJAiAfwC
dTVbI6MfJP+EqY8fJqdrWaWppIrI6EPUOiqMzGL17GbIFZcXiWXA6jzzNqIm2z3jLXBYsqKrukM1
vl3hasJZUkJejKkfVxF0me5AA161D2mJt4VXwPSs/rBbDDqg/573cZu0b9EerKpvGG1EVdI7QfRD
09sldiDBCoX2iYvXhmi6003OM0w/3u0NloznAqZXjzopBYIU/X7a1AU3/5u0K94x0o/Yg22UHltk
8x2KiXcyk2/caac8oM3qwfFnyoFRuUK6IxBJaI9vUwAy87RP+5kbx/eXZOI+vkzKJMyPqrffDNfn
OtzFpTjcTGFv+3g6Vf4/X89lHN5YSLGOdQsd+jIg/c5FWAJTviV91zwxyVm9VDTO+dDfsj+kRm//
OoCPrsc6444fUZpeua6+vFu/YY3iIEQJlkyni4Lp97F/ROfAJrC0l0N63ZxJX64gqkLl7sI1BKY6
FlM4dSiMeTYisutlol1zpnvdA75KJdLD/04ZPkZylV/i9Bkbbj8nVIcbu2DJOp5fu8L8Vuhd4MGl
TnhQ0ODF1hnee99UnEJt6iTicx3Ry8jamHObTRBJHVEDmNA6NGGCIIhwWP1YsFbph/9HjgIqSVBA
e5SjFbiHxtc+kuaXUwRIHLhus37J1Sb79wqkUDSEWWcoztGOaAwr2OMIWfyypueJ/gkEQoeCrJVp
iOxrzTdKLYYDhN8ItQWA5vR2wZ9hnZ5e/Zm56xZzaEp9bKSoYZpEHNJKcaovsd0QZ7+WmKKgPPrt
fdJWdQyeGhWmU1944244O6VygJ35CblJ5kJ8otCskKRqUX01GMrqNydJiiWJZz0EklzsIFseHNdw
LOeyi7wV/AjDlwSNERZgGe8Yh1U82wiTmH7JN5qnDN9Zfi43kUm46d8VGYiWARut3mqvAyKuK4xR
MkJ2lnnh+WhjVscTkHtAnMfJpItAgMBo4yftHMOFqsfcQ/FRO3mmKhriFlrhc2Qy9fTnqFJVCKSi
vEDIRsJyWuL5mNsDKTBdST3JmICzn8V0le5P86rt8nRjVQKZUr8UGCp+/x706e/PYz42u9q/irpL
r8mDkDvEcuAWY4Yv3+YLNOba04UjF/jZu9PpgSPUUpSnIpIWuH2uL+8LUpaV9AJufOArM+VkObfx
Gf/Cr7UjKMjhXLgu8B3fjN6uS3pvpmpEj/TiNIKFOpNaXe3iOtZWPOz9hlAuojgXQpOcHRmFEKRp
FmfiNVVwj8LccpLxYl+IVqMx6kxRcjJ5NDT7eza0MxAtvOMlkcbeO5j3ImH8OwobQsEI0UY9L0C+
dMHANmMarLhodU9Q9TkjewvovpyyKtHGTNQC49QFZmb/TK/FBSQ4aNfDLZ/j8EK9qazJ7P9vUg1f
noE75qlApIqAnC1uQ+jTfs6kKPvd6YIkl8BJF0NTboueqttAtFiEisXDvXbLIT3Avfh+HGVR6J3C
Vpx7UfnpSxkFRLBgTcv/29KuQkEAo/SFU3RtYquz1e4lN2yGeJGSaXUJnhSaEM2YqED2KvkwS/0G
q1vUFBCRHwJ/bj71ZM2L41hhd4Xr4ZrxouK1CO1cNpBaUjQ7C3gJkpEM9AopyjiJ4UcRt50FAm9/
PMBcUSxoTD79bqXJ+TgeDgMgMmcA6cygBQTHr1tochE22PX7HrRDdP66Av5xnFffCbIa83H2lfEP
F08hxqQeOYWksvl8FIa0bd+bFH/aYAp0kkIuauMyJP+OJCYRKnHZHD/8E6YTC+coTvr1Kos7reBd
VbDK7AoAoYJDG5mR9H3G7zhmaaGFHOuomq5q5G/Uvt2z++U4Mwlg8RHf4TqIyWKLogm8rm/eEW5Z
8EvyjNpP35I0WL1mPjxtGIhVT2oJXjdgDdrwp9jkyQE85OMaymJPusLu9XtCoKLwZfcO37VJ8CZA
yuNtYtY/G3myvPKZh+N+/Mx2Hzejg68nh/jiy0X9GstqoumSeu1xkBRY18KBmtooV0bJg/mq1S/Z
Gu1K4ap7METHbCC3LEQCEorGVsoMSvUW7xrm+ar+1qAn2O/4y1b4e7jJwU+/v0cUB31ZOOYhSGyI
sT0DnX5uYfBeM5lUofD7QdnVpKt9759rbi+Wv1jUgYVyoC8cPEakEcViPRLJEV5Pxk7eKd+9Ne+b
ZeLFtWBXNhnVyakvxhVtyrPLIbzOsmiO3DGq75s7+El0Qyq0AX8pZ2++Gl+SlUE7aqa2ifCaxKO9
Li7JQ7tjSSwTeXpm55NaTzlW1PgKVxqFzuF8V++7hyfZmNFHfGSmQNii9AkSY8fJCzlVKO3qVFML
1J/2eVwek71iMoMyW3VU2BAr6b+8EtgV3NEVw8LZ2edBR0BiKkq2PWIWKA3SMKyTeDiERBmOuN35
jI7yoNjbzpEaJJx3jD23itkebpjIHPOzk0d8KQG9a2RpyzNhHT7dfJvq+YtK41IbcmjxEayf+E4V
tEMwqgYPBONjP5A6K0KInfvzW9oMwD3rzofwtTnKYtMnxLNUPct+qPnhQfPKQm3GrbXouuHRSthV
zimkP5SeSkT4PqS/R7B45YBjfbpwh/m8CBec/HGuBCoCBGoIMiT9TgyJPCE/WEkg2jX1ZBau/IVX
k7ElSJmGREMzyl0YkyRSYUmvFqN7YERI+srU6RCi8K1gxtWP3Udbgvk/wxpD9gwLTkEYunpilh7j
AsFLa7RJzQZ/sGuas2eBEZb/cuL6eeWUP8Z6Rwt9HzKErksIEiw71ZWPuJlcr0rGSjXniz18P/QP
sm1Qdr4DdcZDAN+dz04UFWXAQBN6Pb5GolF/2x4dzJNPToB7UZTPAJaFXG/s0hIjESYVNMxpjvF9
TB6w/sLnFQZglAaco4mzQETRMc3eE7P+CegyXH/uWcykL525RLapKARP3Tpu6QabBSVoAwGLc/q2
ri41qhg/R6q2nJ3sd9iQGtNeSSzn8YmuEtw5t8x+NRxgZZTO/m9uf2xO+uuyTJMs9gzd7FhDG+n+
kHWTq7n3IhyE55dksepCqb3W+320+zeh8zo1eev36mvKgvLCWdfhMxy5HzvX0tXYQ6YtxjKXAcEz
2t/8kPmSg4SE7nfs9k1ezYyeU85fuzx8Z/3Fel99niTCT2a4BJwwa4CQ/1EfIG+YCfNTplhVugCB
6MsHmakuvs6hlOSQz3g1WIe3PY4RDIND40VeNP/v0FUAH3OfgzM7TZe2jal/yO3/mjaMOqMlxzN5
ZrwpyZkQMLL43rWO9NiiBtmvbDBya8JQ/iARXXnNBGlLXcl1F2v4BI//oeICiBx9laWR74R36sIf
m9m3VIx2GGI0y7c7kAO9bxmHqGyq2AM7Rk8bF3L1yQ9/BSqUN4v7Ukt4F550hr7p/cBxAdLieZg5
nGermbnZcyO1GaJGzzVBjsN8rFGDSSzDm9+LCNKZtc9KRG8tM1NObEZhRsQgDDVEqXZaNoGL0akD
6HgSNN14/Of6BA5P3hJn5Ji+E98yyi4MeTnKhObje08Fkx6zO4BYAInaGspLQKuxBeCBAG5bLb9L
VSwaWG6ujAP4uOM/OOUEee8l0tw0kqp+vSFSbJMvxmbhCL+w5ggCHuHcE8Nfn54GDb2oT5vxiEIq
kHcIDaMVEI0jEPEjECCVTSnSsAthi1DFtEU+6FAdfVA6AZLpmJaLxzcEkA5WqHPIA+fUurOktw9x
GAjrLAe7GqYYAUI5LXeZZDzjKoek8pnlgMUnEVPS8bIu5Ju7WvfZjXwFS6sm1U8GAF7qTS3iMUfM
5MYEUlEuCmdkc06m+YkKLnxxBGpcX5uoDlRLPNkAQrZ4XjP5wdyf9L++jRkLaVYnOa/W/YWkgwz3
3Wt3gaUL+VK2IRibu4tMLMNHASChrWMgNECqxNQlR4xy7NXpDhCH+k0hSCv0V08X4A7J5UPNAPZ/
kClmksrX9OnVHZL50ZDHAbenSXKS3RW+7x00D6sSCoV2F+qgOnbtIbcZPeh/+ppeMl8AGoV5RDNh
zExvkFL/+O6jngpHE+i7uWZXeAQYSE/PUndSuX1wJkTJ4VMN1O+qxHMLlY+EKilLMkcMBJVNE/pn
/l9nrp8Y9Vo5iPgtPUI0iWUdQZoo2F/LnPDEysAi6t0Uqws5XTt2i818VdgFTQ1lDwBfxYnYvyNa
FQvhLJDvhqoqdx2IEu0isN3xNu+kTSPWdNNxAioDdnS+IAl8nrXVsHdoXCiBufr+lcElKURSKKZm
9Qg6zN/t1122/Mdz2bLi3ARHxlJFTnYVlPq8eJqM5jXHNf/GuX6W+eZE9U4ah62+tNt9nwNGEB7O
3kW50Iy5MGLwS2OgqR+Nz9iUwphAXKgrMETuEf9QN97n4zbv46nAdE5MeoIZGvcMtIqkleE13zFd
sNA+dXrjz8OxYPMwq2+ZjwWCsHeF9mp2Ok5X43GYuvAlQl6cWcWnaCEgxosu7nyIyW5tuYDsY/nm
zi2r3SBUWYbMTyLAxFYYogX2GHb/6Qfb3nLoBXvpGMr1MYFkKw6UzrplsAeB7MsoUdFzvb+B6/ut
IXkZM6CVW3u7s9wqW8F9sUJloAdYptnfDjHOvBqqz5OiUDWq5uuRwlJfqgPgqGyySjM71sWQmeWx
p1xhKBWZFyes+EWXkUdB90hGulNavEEKfSljdCaJ/+qBHVLBbLUHRft9M2oznV8ihSzg7pr8a+HV
xJ7GUhaciXl3o4zz7n9mXT2a19EMDRJ2CFCK4Zu1U7rPOYl13M6VJv9Z1epWs7H0RS3ZnWujswl2
1OLxhEe4tmO1W5QuZ/Q6gsZlKJ74Ll2h5sgIVar6f2ZJAtr1BWB9oUubYUrjOfVb/dZGChUwumwM
1QwNab0nYBLw4AA329AGcHyKFMV3Ob0wSmU+CwJcgNJRDAC4SQIe2A0d7HKNUq6v6SXibM9lhNYP
8/S2RbU/JhuUa+6rNw5BJdaC/u0bpvpenoV6nNZY+RMkgYK7BgZB8ACZsll8qpk9Pjju7ZCJn5t2
ZdbqjFuVHcJqJk4KHyQ7AxGBcbfXshQysJtR1XiH22dMxSndjPpkacqr+2UClP7O7QyRRjfD/VaG
eTpHLmDkMes9oRiZwLuAe4QgeGI1zajWww+f5SPyhR3kVDpU9dSUoLe4uKpe4GRY17rLY41qu78W
77UP+RqLcWjk9EG1YRXzYoK9Eb65ftrrDidl31PZyhuftOep6euiGcHVHRInH4tVrGt3HUm/yq3h
qHL2v/YHMIxh3FjtAxB5wrvbgnA5BfxSeu1SjSw6lrDApdSzg/axYKUk6JH1i2x/jPuL7utui88F
aD9hx/YMFEE1PSDzDAYI+Lzp4ktuy936W3pZIUw0p92SQyFNOmZvx2GZPj4x1EhyZKh4gxkaZDyb
7ZgQghDeWGyhKSCrtjRrOh1SCnyazvd712dswz2DsNuMrcjuQDrl9hTmTHtof/GuSnvZeLnvTaq7
W2QO8vip9stQGP9c5r6TnoVTUlJzjr41jquqCY5BBvFJLJgLx/7CdpAlYP7MFWE4VpA2kBlvcsAG
Hn5JeSiz9RSRtwAGO5nrroMjQ+GQZulFglz4auDYW0yJDGtqXmOVL5PE0YcnQxDhWmXTtuR2GSeb
HaJ0w12k43MJYD/F7LmD8P+Fdg0Ojh5QDGef4uw8ZPcKR6pFqlyjyPJIvbbZZb64r64uKnDhiQV+
EUZ/2fVfovgTuNjFalmX8nHci0x3t6jU4Qicc4vdONN+fD0T+A6PUsvmCT7LG2bFw7agCwZAgim9
DtK8BxzDul0XU9Lbe76VpcyYmO9hJO0ft/aE+AgKIeUNimBXmi1EWoh6nBzWMi4tYc+qMsIMWo3P
03LyOXJPjpB2YAHg5iNzuxp/jzPuKnap+dADt7yFSZKyhottT8Mb/FbDAS5W6ZN1qbEhQn5FzsIn
mAkzMrpWKmlDFEwMyakC6z0Hr7cAdfe5js5ACUl9d6YWK+30wk3rI2Zi+NPfAHRxignrl/YPoaEi
TqC/SCRcPDyNHf9za9mWKtshbMC0NDSGxaSwjfgZl+pQrtMDHZhOHooEKytCn1DhCsQihUruclT9
PKOVg5AkaGA/3wZIxstx1vd22L6gplEI/e9LG1MnFWzCb6LLQGD6ssvhgBcHQge7xqJV8yltKh2x
t2AG1cs2MTjU2eyRmBt2vDCoErYyHG5ZBgF/4oBUmM6TCBj+J1d9EU0kyLIiA5LMCU4IIaPbU0Qi
ld+/WigxTs2U2VUlOmUwXJsUdz9KOeGJ8QsNl9HHa6LtGSv7iWSeo+yMqMjVqLLp8MIrvTF+gptD
uMwi1VAmw92lsH/n8Vy1+J6y0aXpJGuyKdVdn3+Btt+JrN1iwCQjmnlU5aF9yBry1QAu5vetwkFg
SPYlBRw8ItUzrpqmz4ecNic6dLLIQgqnw23+PObYTEznSk++MAyl0+GrN8N4R6AnniCJDgEM7ES1
ZX9MfytLDJMvyMTYuMx6deQbDyyqGEXbG7V4lBFRPDrk7fWQMPFw+QlJkzObfyAVqOOAHYsEM/BD
EemJBI5mwNDTHqWNvPOilbiSrDZDjq0VQHSzlX3a5gXbonSg/M8ZoCDXjNb6NjjKmYzwiGlxMGUj
EYjmcJahAIe4s7+YvWAz7y9mMBTBvqt5fOnhEepR6MZcNNfSRuw50Z1EzBE6PsgoxcwIN5xvv7+T
xssh+MxuEmgcOZA720POEgbyDO1cW3n6ozkaMcz1LeWvLfOhvMBSQtzD+Ms2gH59W7OHYshr6NvK
VH7BQR4LBG43go3SIbpmJPj/KPLROmHURivwg66z+ovcbagsNGnHVTC0g7xs23jJoeIN+bBkA8/c
7zMDPkEyH1QeD9QuyF/ils0O9cq28tpIE9wnuSGGljKp9QwDWcaENsA3IxMBsV/FLuAE3l/B1lYU
RN6Bz7qXsRU4ZhqHsa5WAau7TcJ8d+YRiBDxQThPz+FpCsYtt7Z5FYbu/I2MrA+/K8CbGpYoD+HS
wXMtWMmaRgv6HVzVO0nhKUFxpW0LxXiLWNCU4NXrcHhhFvPlri/SNL+Y7DU282eP+OzquFaDxpOR
fxPPUVISDiDiGdlGdy6sn5Eo/LhXXKhT74/CiknGsJkSHVDKLex7DCXJSWCkhl+Eg4UyUsFtP7FQ
+P4x//sC8FIFvo4WQrZ6MZMTUMpUgupqxsMV+umnGhlfB7txC7y6JuaLI9uZj7IvOvFnLv/H6Dar
FcM7RAqxB+ByJmuz6+D1sXtmPbb7Cxhv1QpBi3wKYVlOpo0xe91NYgo5jm+ZWb1sWX/MFsSt3lx3
byRyR4OtAGl685a90wckka60mmCigQZyPumHxn+nkZESyZRilrtmkNcP0cGS8IGxaUvoUnJUwZGI
BkN8PMNO6gKXKFclQbBh7LAb+DK6oycYxOqMR/aK4KkWIKZC/XExu5jvE6uifMQvJHmpIrbLSL8U
A5E8acUwFXHLEitHSEdxLc1kn39GUHi8klH9QxVPw2WZRxdd94AOyEfkoGFIaF7ijv9D2hmbN7kf
mjBoWJI3qxs8GOZo9e8S40jw45tFIrcAPxpabKZuOa4f19pu2WqNf3T/5lehSqvI9shGhRctTw7j
SIVy2B+T5Pih25miZ2nzMygMYHnNlP78kWiPsLZLfS2g9gy1Ser/knkrTnZshS8H/Q3T9LEhh0T/
ljvMKlbDY5JD6JIaODbN+UKW7uUdJu/c0tMKi3y4lCr49/+TK+atsRQIggxxdMY47WvSgXJW5URG
7ah3Zh+YdIcCqNCVvP4g0BQQcWxbG+TAm7SfJ7G3Y+rQtzRLDBN/B42Cm6dOdcadI47QsXwAyiLZ
pWL6cAaBdqSoksAGPZLE2HJ23ENytVm/D7oPiyZN3UzM8gofLjpqjN8+TCgQmgaZR14bZaesPbPP
7kZ2Yy6VHPlC4zlBmAY2kTrh0yv9IzIr8w1UaD9RFSux0S33wwuQGm9dRZbw4Mda2vblKeMNm6Nw
GAEFprhy3uStzac6xTaLY8kMIs4KS98/HCjJvmFEtqqaTG9hGdP9qOHEZRlCGXbwGVyaQObPDZfm
IO+BuuWQMX3y4gmVl6u5qOb+Owo2CFFe/bJR5PJhNSgo6cx3N95n2oFlF40vEH0QTFc7hE9pKHwU
BelwpbO7a2gQPH2RjXyz73CDNey0jMwrq6F0g+XLUduwRprLayEOlsFQej82LYnVe0ckMBn7gq9r
a9ENdspCtvqMGMuLWTXpLDxVaq3e9L3vBI3PYYST3H8SQGn2F/Pb0vGcz/QqgXqGKgdyAC53h0bs
Ca2pDbUAuKqJLiK/3rzJSoDkUoUgqlCvQQeKaFwjdQ4KGmh9IXXdIqfx5IbVPhWPFcMuH+JqGBuB
vOojg27moMB6GYKHelicRRqCtdfxR5S+ocP87lyoyewjXK3QZCkUQJz2N4ZFQJsQdHrL1HyG/yRD
5920emxgEzwE0gWpGbs0HzZk1jGdepug54fRNKZzaRNEwEQbPxvPR06hA9FF10IFbb2L+EgtikQL
ko9FrI/98V+CRKRUMydJ/2/dhvqz3JLzVD0IVjth4tFn88ZyLsN2xwAouTrLGdT15n8hZAV8lq+A
zgiu111X6vRGn++Iws0Xft4FJFfVrmLwb+Pgjzx3LDtirJsYKEOUwAj/uiTquFCzkzFda0mTqhdN
rEPGyb5sjSW7w4mxuaPrR3PuZ+85bBN13+RwotQOltxxKg242ZVBSiIIPE/blBom4T5ZOYbIiXnR
rJY8zU/0+tTEnVPLbh0HU7QE3fX0ulhsXHuJSQNgoIth1bCCyfbkmZF3Kzsj6mnrsB3l1lYOM0Yz
iE86sO38KZqbIdzyQYu4jV1Tbt4+G2iULPQSVgfmxnQI5Kb/IJm0mJ7naPpYdp6LQxPlo/0t+k0u
gUy3Kx5gxU5iPbO30kSrkQR6SIscQ/lkhPmCK3xCnxH0yh7E0AJXlBp/gOPi2XiArj5ipDGiDnAB
tBai+Fid9opkm73qIwNdgYO0Nfa0xiS1PndJusnnIXJsd1qXhHB0AR0o813TeZDsJC0ehuD/ROcB
rsyI4H+K/wAUX1rR/FHanKYHEmuAyuc44srDQJp/FhBM72j5wbmcBqTRAQZaNHcpZ6N4qyPLkoh4
sBV7HzXtOBCt59xTkafMJFcg+f6RJlkhZlceuDHb9RoWakecmwxohCOUxflA0XMAUWgPusgsfHBQ
i4uX8EHsHw4y5HlcsbPBOMEk/10OPcaSpVLAao7yvC6B2wn2TaOTZoYOE0snlZd+VsaevHzvZ046
7dU+3gC5fHPuoOIO/yKQ+5JKPQYL3/mTYDrMBd6JHaHO7hivjoVvEITFGdPm0Wu0Z86g08zDtnKI
MqYVMPjleQNe6h0biIJCLBAWnEMD72+fmbZiGGFdtl+OnA+Hl6iziyT3t6hj8hvxhyRooLLNEyj8
ZALqz8sSgzo07Ks/+/4lbJfW39mu16Vgybk8DxDduSv3duUcHQ/Bg5UutYVADmwvdaSSUn8y+3Wk
MWWBl6ZgkTgbgrqwzZKTYPdEJw8H9EqnMJDIv3OCNCB7hVTZq01kS2kV0ydq/PoHqNZox92qoiNI
UrgJ2XgG1TeQH1zRfLBuF/zB0t/vet+u3ei0zWr4Rj6AxeewOFiZWgsSSne6eloT70iukK1U0GZz
ZDfGt7qHvMqcAH057vHhG5r35xG2OFYNggF3L+W4hWfVuwuRlgOtKU5x9YbCghbCsZTlZxDRZwSi
eMFJhrxUbtTEtun0hGRFbblu0Ue/dRMBfuPf9tJb6MWP4GXdvLCgAujmAsfUNR+2lV4nCgeZxx9M
H878GJbwPxzW1G6pcWy9TL8ntiKqVfaUdh8sfuSa/Me64aZHBsRIBj4RDRIlnXsfFSPraNPv0m4E
MjICoWF3K6Wo9DWt6ZSBBWH3L9tRL8Ncb/u9cbfpFUKAJH1aBIqTNTQ6LI3q5/hTKx5FTWUWqQrk
/hZPkP+aLVYPKBNdGQMX6tkPZJe5wJRedze+EmEiOedwiHi2qbvLjVd7j5aZmwm14x0VJ8IQkeh8
bLqW85aQjCSikcRaEnEhYBiABPTgUQnGIzP4yLAUqS34EEeYTpFXuHXOkRNA9WukUtVVP6FfXzO8
MZAdrJgr55c5p8wnCJHZRQbEQ1qdKRj4VwKjwyMU2URxA2+64XJpkW98AII0rnAG/C0+wV4QSCON
omiHGZsXi+gs3vs8elIXDOKucYTekpXrucC2smp7qjZ1h93YxiDrdH96Z5Xd7BgrEhisvQo2JG0c
F0zbwG3VnVXf8lNrTnpfdHhEZ6Av7YNbVatQUwIW47mqHuB/f8MgzbMeYATFssH7VyRoMVulBhsN
2VdYIYCwA0Wug4/bkAFa5eEYcXVaBqV7GM5VzQWZh7i+ycqMXsrFCyLsbrvXHLEO1k53/At1jb97
xSnSTrwIh9qxJc2ZHa1TYH5pWeRFAIxzO3bFQWWSulHJrf4HScTX9qdcX7rV7MQgqqezv6P2qAAL
CxaVAdWnMO3jAqy1rzTPKjSj0AnQo1lxuwSk91KQBpRvxGIfzp97f0BL1C+Oow3esyw36/dIAS5W
5Z7hGs5Ujg68RZO62aQUtBTiMpbgfAnv/cjLP4+Nqdk+6xuLswIR4uFVfiplV097rsgyQfeU+D7C
3KpJC/wtRkaSLzpyTZRwnj4YDo/+AmX62MMRfOgL47QZ8cTJzmbkbthEE/pyakUx2s87ykIqwW4v
GPL/pQBfZxP63DIDAddrLJtrLXra2lTaCWHmxqQkRmpHJHrFa48TM/RaUe69kByG7X1qWQFZEqmb
Ya6mxP6cY9EVkihMIudezsBbKEO7r2H0OxYG0nnh0ss73pdmT1bjIBSRrmCo4bHOKUeyaJXSaXG3
URponuR6NITayLA8AY3+tViNODGoe1KKhnmaVgc4UM3LX2nVDto3SS6rlRarjMTWAer0V1cYOmVm
jZEglVFnKGcz92y1eKU2rFUgD4wD4Lp3bADBUWcMs79IeMS0MZgIv106bDM4/QQpk3ceIywgtzY+
R86XKG4NmTdlvfobV7F/bXFURB4E4EnTKFPLJ0wnFylcNXz67DT3DV4/pGQmEFlXK+gUacKhivtP
o4/sKn0GeY7BVfacJ8EwmqWM7H6hABzM9RfZTDutAoQ+SHyTNuaDp9pd9rfn/k/mw77mvQjy80qa
4iJ05KK+0fx+/NUg4AiBZY7alJFUsksaH4Vjhq+veKtzfcXRga9caF6aj2GRYo8zFRib1h3mDHrM
8Hqo2e0t0opk2pQACsNThcofmqBGf10kJk19N6R9POOuoBFDvPGKJH/JLWOYhyS2irFBHReq9Ev6
TZXKa6EAc3QlrRu3bRjBQYP3wi+ptLEyHmIRIRT1C3MxLZB3Cqi9hqP01FoMf8Iu+G1Nb2oT9IyH
WuwHyKr6ScIk++Lm2xRNI04YIuTmq8QLMQf0twU11DK2HRVaBc6OGeAkDT4V+evrQ683ilwKHNDq
Fm++v90h3Cc3xrZk9VsLhHKjzZHvZhEAbCUKsfZS4QKIi+S3fma0KsY5LjixQQjEeX3WuUTVJenu
WrY10Vb3R1eoQ5jLqUDzcLeN4rUVRFvv7KmXUpW4Z3pHX6aGBpw2MzjFmgdtZUmnUR1wm6sEkyHG
suBHBWpfcwTkh6pBe1w7/PS4nhD6fFEdQ5BlhBvJCI6iMjiBz03fHep6h2TC2OkgHSrjVga30b9v
s1/V7n2TIpLik/U2r+g/snX8shqaUJrbnz1OuO1epnkwkXBoWkqHVYOwZ1WiSqw8fxUbXFgJleXU
IfNTXhuvSk9dbJjnRLZwd70qlbyuk9Hn0q+lXjsD3omiBdriusCY+0NTu2mygFN9sqFSGKjqcpPW
ZLrRiJ5MvtP0U/o+XABjltCTijU7eVNhtpwqj6oV4aWy+L9U8WsOsjTRYoff7QgTLzfUIxIzbI0q
Ct3CpEI4yVcY13e/Xl0795+sX7N9kRwR4I54Vnv+UiNeCpHz+SO5+sSLMDOWrNxA/KDZcWx95Euo
bGG2p5B1RV8XQjypbwDCQYi3Tc3qA5lJ3/SSP0V2CMT8sJozfvcuKb0uk2DZNeBUG/GJp4a3hB7I
4STBy5o5adhmL/df9zrBFymCM0+l3T/CD/3AK0R4yBbz0FUoS4s1OKEWL11G6i5wFRuueEj3qS5j
a9Fn1If5p5xLJmYC+DBXwPwErklT837dSGystin33VzBNHQ2z85R6QFjjKhEDrt5FlTOmXWyEOs5
tfi+LV14uJaQzpPSOzxp1z7isagoB7JXmLuAEXlMcmQbNc5cGVotOqajditWxPlyzHp9O/ORr6+M
bHjNpW3Ylt2OYSjSCoqj0sevnPeG3oUW0QXccrEU8F8cGYeP6ZXHTE0p8k6+Bo1jmCgDssPalrcy
/itGKESFhIipYt8VkUVaDw3oRnx/ZUfHZ5Dv4nG1Z47e7ToPePqrIKbpo8kG0yV6s5IT/2jfe/Po
XzvKXgtQ54XlJZeEMo1xE/6/Csslkf+jPYbXA+TjYNPqdih9IytS7pbbdQ9rNZmLxzybtKRDSBfx
QSDHGv50ki/aZnDjUrAXM2Xo+UKw/gnVCyJQzxewF0bq2lyG3yGZDncbkllKr87QTzJem53gRqLP
AiRo9Tv5JTcP3QXbADrrOhJIq+iUHvFYzgcL0yLxIvSh54ORac6ohsOZMBq0vKPy9yJ8dBAvN5cm
iXTjqDA1XU7kfH8NkgMULJvp7FGwHzKSkmmwGLCc0Hv+L4Rc61pez2xTCdvwu9/Vp5jefllGu65F
XGjtJXrmmfgZOg2wqfwWIjlgiBwqirNKW7CxlU9ZvFFpKblIZoKoYmU5flElu8YDLWleIgPMf7Sa
qrNbAtBeifhV/iFfq+ufeMkjPwN0aYPUvRop2kgng1K0+49uJ0FlglnNXk+4JiemJiPzPHnRYGZP
kwNTOKMDBWJ6Q6wsbxEhys/YSdgejwIu8sPkmfWkfr45l36E/rwcZ16cMCFlUdDbp3XXY9FRYaqf
xyY0fgy6C9rV7xtC/6iWY49AxvqRigPHFuFrUyG1OJTy4FsXylpSkQizOiK64UbgK05rjdO7iHFn
uHKHSqUjxuC4OaoOQNVKr0W9KLHBI8dKDPydvdavD05zdAY9zb2jHf3hFLjMit3KOaJlQ8MFqKIc
98XTcQtluoWckN+B2C+ARS25H260lhSiG082YgpN6lB4xEtii6KSWDeohG4iv/FaOjZr1eOL/vAP
tMdsVJjZVWXDWNcK8fnzIgMp7DY9hISahxIO5x2NEQqXRWb1y5q11HtXbQlAS4zCv6TD7o7v8msO
91DqWjwdZKJY7RAK83i9Svrw9ToabtYYGIDS77OGsTI+4Ux9F+zQucin8WFwH46tvKkhMcRAvIhu
QOPE8pUcml4OLxo3CN+r+KW7wNMIxW5xeUSvmL+XMpvAwK+PygNBQpd9Az4tHo/uQY1g9U1wZYk3
18rUsPtVnxlDS6p/UEhq3JbdeIl4WlxQVswOIn5/0U92Mpmcjfa1wH2QYYKYvz27A8Gq0g467CrJ
ElXabYftQS5662qnFKdfc64nHphDo6/ePx5VGHCc9vuiH3nZDqe/5+4FkGT8XQvdVtZa1fJyRBfi
VeVBXlSH/9p2tSgzT6xJkTXqC7n90OZ2VozPzekTQOW7qsP+PwqObpjsGPyl1vN3FduMsE+YhLly
LTAupukNbCs4HrfUH/7RUx+t7QuxcdJbJ2kDlcB3cSDsS6gYKtFlLU6kNPVwUsNicePFyMG0QF4/
ABnv3vduy6vA/8JyCsKkR19nDwXIrZ4m/KQ3T9bCbuKDhwxXBpyR9Zt/JBg1XoIash/fteeAV624
PFkln7JNXEDYciVL0GkS2hQKcjo3YQcrCNxWG7b+IhE3fEEYYmB8m3S7UJn4eS9WUn+OsFXsX1eS
S6Sdsj7wweU0h3fmPsqDxtAupmnJuFqaYhEtEjNbAcK6xGHBjYGcQUEEaD8Nop1pru64HZbrn7K3
NpK5qNMFa0bBlo5iGRz/YM1VOfY4Sa2GiouBHA2dMv6EJmuubxjM9tx4CTRLNZGaVU3dhp1Ck8Uq
lf/Bwq9l0TgTOriH8ITifrmLiSKx3W/UHGwVm265Dp3FRkr33dAVbQf8dxotIo1K28MPvFSRbwYK
Ea9aiyM/o/oBtYkM3mJB1Z97i1NnnZxGpQMq2lEkV4bxGdcitYwvwRRxdEhf7dbIzZO+nU45Sv7g
Su6xTx+UDAzfb/sMqEUDZVbAmDZO1xM9pBKFScIDWzO6z5e5jcdOghJlPxKgpX2AniNqg1jTi9ac
WIc8vvwskmvxwYaApRqznt/tevmJtNrL7YbVyrXsJkGSIe+Bb7DiCaCxnF6t7JcmvQ3w9pOAN4qD
+q5ADl5OL90RTHZtDa0jyTHMqpfKHT1KGJo0OuQzMDg8xwexYOAaI9u84qbLlFn/IjaSDCOwloqZ
2ohxGyw3iZTMlMcy0tdkzoGuTXFYDK/OP3H7xg+drd5SOhv4GPmOJnM0ZjLwlQhumto3cIcEfi5f
yha6J0i1lIgmvE4k9JmF8MhG3wRCtqqNjzdWUzPbQvWy0SbR21ywJiHVCeZTqiGoh+ltc+rFsNJU
7Dm5GoXsrSgzWUFMFN5/a7sWLztVeajnOR9s8ccgqcmfLcvQlU6rLCtHQutSSg+zacM6CyM7/Uf0
4o789TJoruFQl+ksw5dn/hHFsLjN+pspJ+seTskdT/REKnjdYQz4Nt7v4/69C8ooK/a0PWt99GMQ
yRoBmkjpfn4DHGZEMaCApf2y8JvdWUazer/22wUqWO6Nz3RKWgaOJtMaHIDC1trradlrMLFNa+Xd
JFB4k6SUMCd0IFyEt1eBjSlX3xmjesKO8oRoJceVZm0s18W8728OpR88eTPGFkia+bz8+pEXQqGs
sfoR2MMAtX46UgtHyVA2Q+MPlKBiK55xPLRihJLOdGTqFgLumiRhFnPC1M5CRWMFH7BnOLJEejdo
tIwId/HhqK11hrgRG8kfpdID4cx9eU44QMH7c8nhHcdw6TusBh/YvdF61kuCH3akYpuwlLIWilnd
WD4OWCdHSPOMhY/Lwums0JP8r5feVf3BS8UL9Or8XUytOxoGioZ8Y+EfvBft4re0Fk5R5NW+/aez
D3/Y/MyCgfAFaWkyXb1HM/VrVKlfu3Qx72NPsI89isaR0/wPzLmfddlZ8cgiKzBs+Jh06qoYNcsy
PibGjYRINRiLwVcWL7RGVgYjq6+OzuiOsRufz6WI2HjJDaYeTTn3ID7soOSd5By0pVaD4M5K6Nh0
8nDSIQkyWNJ+kOl5wl+Qo/pTDp+gGR28gSl4Q1O0EDTT7L4oz6fbtgu4cjZbzL6dPdUezLzZAITq
/ZauU6Bl+Pdt3E2riQ4loPgdJSKH7l20TWcbilSKAL9BM+f+cT+3D+z1Y+RGVFS+cRqQBn8uTd0s
JkB+aJlmmRM8G0nhfF1ByVzOIC6HorPsSef52LCLXmX7x9xMjYs9oo81UGhwA2ZSaXoG/K+IkbZy
QPyLTIoggNp1WkRyDvCpii5buB4LXju1W0XEfiTmch+g/XUlg2d/PSwOAhapbfQrwN8rK4ZXuDAN
vYiGYXk+bKsaZUDCInwLrfAszwVPwmQn7W1Wgy3QXK8YFZDCHI08dAfk7nKwlPZz0T0BJq9oDQ/I
UazEpKqqSl41wKhZL6p+zF1Uwc96bsa7d57RJBbMhjmRtk/+AEwwKw4QXhEZi2XRVc4FTXt0Sk40
Uotsl+tWTKYfpRJWnqIuD/2ZnMC8y9IVf7mC56EikK3I+iQwXojApKk4mDAAc1cceyUTOH5HUo11
+b8AoXldStD3Smi0cOPv6IZY0NfPVT2wsdm/9fBdvFw57pOSbwmU5yQCfqsj//OVfjwzYhWIu14V
JAYaRRcjzLqqu32AmJzaHyA3VF/uxSidJMa164ljuUMuhzrkYpnpXrBwvpgcWRmkHv1afczk96re
IT6b1j5/nfpSZ6xgtHbZDvjKNX4/7imVZZt4g6SKF9VB/eUfS0buQOB+OU0T9hgTO79ABKSnL32I
XOyh4iQiDWBVEDga8LOVmCxzSOZE4/Bntuyh1kMSJj8gIafvuvDt3h+Ct67cOc4S/sGjYdnvLbxR
RrLa8gEBfUvlF23f9l3ejDqJ94qj4LY3DkraHCKbhfdkm4Y+913NwsV7OhtSR5gr2sNIVFyN0BIB
/87tkfAJgEG/JInbgusXHjlDyh0iD7e6K/NfHB1dVVnykGo2yrdtD3UCzkQehxfOzmJjDDKKmxeg
Q6Ma3TYXyTMkSaEdo/oGsVTDeckEIdT8eZF7pHEiJO/uvApwFtmUN47wki1Iy3tf6R6aN3gb6az8
Izz1WZ150uJwxlDusODH6NtVe88Mg7LrsaP9LkbtzJqGNe3qTqZ/NVpdEKltFV0xhEjZBO4d17qn
8abeohfqLOIbiRqh2Hj7Cb0XbV/VjyrVKs3EuwBWamGse+IlA5wNbA/aLDrCbjh7XYWHfZMYECXX
J6YSOV6S6c4ghQUg4F70NHM8O9nZHxgbY74N7G+YzukO6kal7j3IfiBozvMlp193xX7vVONbuSNe
JYgwVVYHHMSl27ftp3A9aJmJcm1dpFDTHW5/RVksobJnC4zRjOCD1uAAmx/E1Mx9ubGGVKGX4Fmh
848VG2AsEA1HNNxJtzRhDNqG1CcpNNjCHpKr0HRrEUAdmhrju/nXNRwyWMTouJrrd5OmPGEw5wVh
uCV7OTZOFHrawcW8ae8An5f4HXP8P7zYVbkiiKsI092GSSpoeVycQwiawX3IkFj6qBnxKxj1zUid
dcJnLwRq74Jpp8bSPxUy0FA5oBOPciTpZZLzRI2UejezJNHrZp8FDYxD8LxvqVmZuUOUttpt2aga
Bbc04QNlIXFk+URN+5lcOgSY+KDDFnv7VpNTRAQbn6L0bxzLCLKWErii415fSbjmVMvJOwqaSeCC
SG0cv/qGHnE/Bho1TTzOoKpo0yTQHL7VSxh2Su/d6jUTJmK6OpTf7j7MrY6ODLx+tl2hiWNjSVF2
mjDn5RfHM0BmyUN3+uoindiYmHdyXlLlSuNJGA15/tx81IhNCr8VLQIS2xXCn+Vg4+GoxWW6NnsP
aJvgNKON/V2Us2uEZqKMQ0pFHkc7NMGi/q/KoVHaRkkvAGJDB5kWZa+yJHq/qMKIxzaA47dsBQiF
w/Ri4qwgpAHDKvi0R5yHWKpaztvAb0PXF1WO75ugbNW8E/6LjOjRLRYVL/R1NNczq7RyxB4gVh6w
VPYO6HdDudud2ZKjGcYkvfwIVEphYYP2AG2keHzzIak+RnjZrvAOOdQv1SbjpGzlg/h6Fthiqlpq
u/rQmSXaVVsoa+k4L6JGJhwJ1Rt/pOfOgICEU87gItjOWiDkvy86jZfji6bCiJbIo8OihCVvcA8h
pj/qVfGXRR/nI61LBLpp5TAf9gjAAb38mvVJM9cg4t5jJPMi6+G+61X3AKhpLtqUsb4jmNfk96hA
Kzo9Ui7bP8CKoR9+NbwKivEBOkl37p0es0sMU6yUnSYGagtGJbmUZHDC6n7dxtikb2lJa9TZ8Hly
T+QGf0jPqUaCQp+e3fCRFv6o2yHAcwiFL4YI55M6OoS9gNTbwnXaloVrdnv4twOG5rOQzInFcob2
OSb9CEVui4rvlvIdW3zlSElojQp2zHAgHzWreLv5OzUWftLY1pp2wLSS5x1D82Na2VIYBlkhmf2K
f1zRXxRtzj/9GAvGnW4GEeVqzae7SqfIUaF/Vd/NsgyWJWfZWIcgSywl9OCadziaVfkEg/chJeDc
ku3tDNy6J36ssRMkP6t4J4MeBo3lOs7jOSnS99VTEP/Q0ZMnbJ431W4LZ+Qj9qVXrl+8tzC+AzPI
zrTZr9b8g9k52VBbYGkjiNfO5kmwG0luB3r18k5jqHzjapMKTv69GSBjpVJT5yE9JLjq5A0tMoPa
unlEaTYzBjA5EPszo6RWXK/IZSXRsjSLE8i81OIRzmdztECwJcDDnPUAQXWNj+0dSaIZQhDg8CUM
TPTJExtafGf1wF9+sVMR7WetGvQZ8QEydpGHAK2xP9I/KH6LmeAEwZVPbR4ayEEDqFShrncDRqYV
qj50fDxqGxeYrIatsjp82qbZHFegxJE6KP4LxOvVmO2iIUczOiMg2naxuYoJMONtdRPP4YoboLxT
2aiuntxgKC8OKPrODHmuGn3oDAD6l/eVr9cCL7FDXXAwLKD23ZNxgWoe2yCdTk+qM8PBRtkvjYEA
vZ/tu4HP4tfNGifKnuWr4dwMIEgkv2mPVm49aIInTA13hgnpLBKUjlRvqh+qif4cLdMAop5bFNFz
WNPylvDvsb83YOri0B6NcYYiswGY6VeFLrmuJJORpm6VXTQkc3HK9CCb1oamSOR6G3hhoilgO3on
VMsOjZ6ioms1xkMdasG02SoSxUMDvHZNZb36ee8FsFYFPAFVDVGkW/gF18rmdBz2OQdfSpOVyuyQ
qbuzwiOk6V8/+lRm1elFKjoQ9xY62rtvVjeYKUM/bfta15/+9HtLayoqKF+LfUscX7z/GyGEZhwi
rmM4LlcAR5ZPsaOXUAwb9nEfJg6nJMvAHncZ7zOq18tSTaDbEvqpa8FqoclK4U1BkmdsTJiH81Ql
WD/EJ+/IQdOGMvXvGsUeOUJmxkp9FQ2KHOKlL7do8aS5GAGGCc5QSqExQdlEDf+AEWqB2hyaSsGe
XEK9f7q4s58bUAHhGxDx+juvfX6bJi2GAg0DMps1SGDxxr/QhwIGDu/Fow5prLGs/LYpR4fGgWWv
1hWu4Q14JGgdCQfw2RprQv8qR1+2gqVzJskCSEPSmrj3I3NoowoRVlg0AuLc0YYP3RUIopSdEDo+
/gOW1aJHgmABaoiLGhINSXnsviurDKpS997s3rqDgoxfSolADkV8jnTcVOIOFy2bSMBfKN3Qx/Fk
SbcoaTdX/ZQ3GwFJFz7NkrbEWOIKll12PgJqaxrnf526W45jR6LOWbl5XaIjq0FsSSwqX0OSKciE
urW7FdWH068UZieO396Rwv2YoLQTIlA5G+MM0XOjY/cjAfksj8/KxVfxqC5l4VIzesZ4mAkoVScZ
aPYa7cWOKH9lEHrk1z945XiKIWqkIGqrbdAhXGxeWCJyhfVnH+gA2eBrumlEiKr3IjY+s2NxpmCQ
zbFyzPRNybvNoleJPKZ/UlrDcrSfhP+Xzc41zwR/0r8MyUwMnwVpeLb8IaAfusvXa9IOkcVijJ2Y
dHEFDQ1WLuJ99vSCAlfJjbWev/phjudrTAkhGEaRbFv4PojQ7RPxUyC93ZXEn1n5m9BIV2uxyCPZ
sj/nd/kG0HgcObpv2nPTRk4G5VtIO5FqkcAKXjiH30z+AK6Zbw5//43jJ6OBoFq8tZDLak5e856m
OS4SIVy3iXrpWjMIyES0DIyVz9O1VsC/cUqCOw4/xaBRBL7e48uvz3MI1eW2fKEich6mE2uqbkq9
D3KgvOqYHNypxCSRrlyk6EG36fvmDWYV8xgcyClLWxslhReA20XjZf71LtKnz/x9lUxpDlbP/mgX
lx1eL95OdbX7uhenVw7DSvzUTDjTzbQaegoUCcJwnS4QMsUPEOF0AHJkGkbTtwdLNlN8O0hv4P4I
p3Nu/sbV2gBkrrLIczO+tnCKlFv9i2IGZR4kmV1qGp5QL2RqJ/xNaCco46uZssj3MlI+UzpzNDgr
YyMzjm9p4uysnGfpBL1xfkjvXTvgNpcGntMhmMl7kmzSCSKyM9HWfp6h/ZnZTxsRgVJpVth8JDds
UvZw6nr3ZxFZpReI8CnijLy79cUWWrDN3BVKU5T++vLjv7gllreVPHswh96g44iB3SBSmNRugPvb
R2fN/5eVQm/HrC9zUN6HqvrVuDuy4/W+kP9TyqItw9yBKChCNCWPrxTIQcokTFgfYgSbE1Lzj/YK
+auwQJka5Zvmt8hzMtzlVXjNqy9vVL5Zm+WUFmgu/fqy6z5JGGUr186C83zJHT+aLTEVZeEye9tq
VgsiRolh51Apne1QsRaS3wvkvA0uBzKN6+cCVlX5vROPRqchpoh7QMRK07JWNIeabe9zYtezEuWz
42Gf+TcCxO87aA5TwofnbMILgfW5Rs43AIeTkdxd+xGiEAB8j9ISAQKiapqtNnIkD3e6x94otTRb
Vbx85ONNn7vA+u1Z0KLdGnzUb5/FUc8ChAhRPtCuDPn4iPx3rel+zlDkoH4fT+lhD2qgHq3EgaYv
2rN63qU7dm6y7x371zKYL0B37MAvXMNtpd0k93XArtFw9THR3jMLCUnQUBrH1DaFeoTTtbqayqKe
fsVWWBq/Kmp1NCbOJMnpAG2IdJEaxhet/ukeEdir6yGw+8sxmn0+n4iUfLjz875hGah56TncjfAy
mjQAvPZ4VOdwSYeuQSTCwRAEuJAB+EtRLxILSfyGI/GlQfGY/kMLgwbBV2DQryAcLU/48PEgMTyA
7e0i6dmnyKNlYFuqQNHiatXkkQV1mjgY3seZAwbXaQThYJ5TtKmc2rkYH93H85+yoapEyfHV8448
hnlNsYqeLcuVibTU5Qi0z1X7df0lf22VN7aDn3qMlp8KLd2JgypYPPFQBv7sMV6p/yqtxymyXYaK
Qe2HP2u5oZKceuwuut37htwVZ2voAX+Kt759htPo6ggHNds6xZF6sYRC0y/kP6999APc9O09Bd96
tE9UTagQZdBNUkfAm9eKQKa/2DYdyALVqkkGyb2OAcEEV6zXgX4+3p4VBA2yr8P20fMU8hltG0jK
Z2QkGAA+kixlsjwshJST+S+5kSF0Islbt9JcCRanblFOwFMCZNXVJqz9Tq6TL7TwrrNHtXq0wvIW
YgJn52MD0EpmzXRJMRTKHjRua3GhiWBhC9AXBrVbpFWN6a5B/gqpmwwb4QojHQAJxmuLikMQrF2N
yoOL31ox/YIDBkANmVqtIUZ+0zCd9zrPqv7vTtze89bihGmDdvwg6F//DwqNX/ucMBvkfIKEY1sa
V27lsrxf9vlXC78NlRAAgZ5tYqCKgLDRsk8xooJlWpknRgiPCHK/ha15cxQ0Uy7ApobdBKP0ZVMt
5uyXLPp+JuQ5DfxdwLTSaaYt7PAs/PmGKAUTkNCt/2ZDYt9mhIMrJYETAYIwScs4pDOUwhLJNMMr
10mBvpK9RfJPWWghQc7fk8jXvSsb27IhX4fO5Z+6a2E91nmeO/SqudkZA9x8GwAA6RfhIeuwZFg4
Fgqt47EDD62AYh+USIMm0fLgPC/aVnoMzllkpPo7MMVmh3Ja4AUm14IgvCKnuzRkb1eISBV5pBTb
CfPxfzR9nscVMmNe90adTbhYpbkiooYqSvcc0LEygjXv75TMLOVtynZjzvdEbwCjeJLTf3d7n3MU
xjjoKs8RKV6X3Qt9kMjaVkat3lH54gufcuZxuzC/Wz25q3Y1Cz6O6M1nIZo1RoLkHu7aANDeXk8B
R5ckxmWnuoWolzlHDbn1Qs2ZhdZl9DQpX1FZRFLKyUyfk1KFp1c+kpM0ObfwHHkPvlKVbLGUVDAv
42i8niKK97zr+gEvp+qQotepf457abaNj29KE+3t8hhAp41Yv6abPYlNpQ+KG7PTjwZS7rFFkC6i
dlALVdu+sYtgS/J4jnLfjtLdfDvxPj7ZTQvf4o5cXUbfOu5tjrwQpuBZVwB/kHAEzSwtrMOIXihb
RmCtWXN2oy0JP70kP5Rx4uX1g/UmXnuyntN3ctZJzx1eHJ67H2hDm9BiHGcrjAYqvF5fuxKo65M1
XB05FslzWl8J9BbfxlUWy7p4cpcf2XYbwfHOOdKtmbseS+lTF6DKXyEfjt7iHR54n+0oY5SoWxum
mb1Acx23x/r9RQQU0ncsVy5sELyCR8GV9hw1wqoKbenzfWpe3AIj7WzFhH2nibnTTog048kOHlEh
FTIvW3mF/GxXHZVl3npphIBQ1bRcgw4NtrKoy63rpD5SxHcZDjOCkVhrdNEgNmac5dfuw00ggIp4
TfXx+MI3yQDE8yMa5SzZzpJeNPKyARMxQCEbvzppyVTVD7pkjFBOERe2stvm+PV3dQKCSGIoDXCt
3wENdmco0ijthOezmFSbaeQnQMWJQ0rVpfbsuxX1t0PMw7KvCp/ECKllEC3FF/oNbDEM+7ugr+l/
Qh+C34es9aMjVgD98YifcaojqkCk/lIJmtSAJJpT1a2uP7Ngi2zRoJlk94nJPAVizbcV598Uk/LS
MhtZM2g0XLMHgYEylOt5ZoMVoH6M0P52LY56z4ps/8Orr7TfslgfCRWyWk01p4t1SoLEUkrsO13H
8ZFiPx1grgS4fddjHFroUen1sEPYo6NNM02eaVQombNYZETO0whbeKU9qTyPizrDHBkm9hvLtk0B
leM/wiGHvtr4ywpPirqC2ieuUMOoyPyCxOkPQ4EYq3OAaPKHcg6uwL0H1KAORCaQwYwf3McilhRQ
cpWIXhLb6mzZJE1QktCjBnBRz/Zmb6DQSV0rnVit2w+fHW2RpHsTpuPTuncqarTstaUzFTKDF/cG
hI8PuNJbFJ/GNEKJfjIDvipZjJvBs0ef27ktX4XSJSbBhACzvEpsYhucypgvrisPSc75Y/w9MEGU
H1PiUelYIl1oQ1ymLUXzXRpmCMEmW35QA6IMp+o90i87QfSE0Z+Eu4cf5L/FYxNIf9i+4EApOc66
1zBteEv1plcke65GY0JZZ7lqfPbq0hnm4bkAuGZJmGHCk6eYY3IyO+pRms5S8KaCq26UpY1fv04+
o6WATJ7d/qHZl6Nqw4BQLohFbgr/D7WZHzf2K0F2cHUEEPTj7dQ7BLxKt+tU67f4jkgqiCpV6HTS
PCwe4kOkzpwsFy0fpno52tn7Wtg53pmO9Qw58M5Bsy3fe+rEPt4IQQG7CK5meJ5SfsVTuYtGtNVa
mWV4SjuKZCXhrK/+PfKQ6PtqTme2sIEfTE7//srkp8Fp0WD8ICiCOJgJ4YyalonIXRanUblPvwTz
sQqMujrExSVA8frY0BIBZ8XPaX2e9ZCw4sQ1UHPirHD4MSVj5f3uch21byNz5lAugXQWGMjeG7Ta
VRqq6tjghBhTx28B3aRj5vNiaRabrb3mQ5upOqWZ2XEF2poGe/MFrijrplrn/AXym0+QpSFx8QVZ
AX9nhhCEIaUaI1MjmuYdy/InqStphFslUvdKZgoSd7BrOlWBKR2K/a+URfakU/yyiSAe5AcL4MA6
EYnCmOeweFKL8TKMxcSqrxOWuGLxe0J6WaJ3E9YVE9N5ZpytU2Sl4WHjkT4LJBX9if9llVruwxWn
alLlKY01N1O9Tq+X2yU/6dFISWpW1BhakfFWTIOBXUhAJKpolPTTyGlOgGZo6rCk5AQ/shCcNR2B
3dxciL3auzwGCcu6rlkN2ytfMf+eFjAa0X8YV/Edf6PxG+O7O0fM+Vg8cj88l1skJxmOKRn9G579
7Hhpqk/fyMZ+31WflMcoGG2c32h0/psg/GjQaS4S+z/XleXsB4bDTU9I6zKX4EIOfoJa3PqXjVyV
Q6Q/g9jvD7dtuI7RFHbIqQ9mCHFMsb2hmEaN7l1GDTxnKkySyi26SaeJtgUfJyyziwd6Y/F2Zz6Y
71zQlZw2QHahFFC2/iHIaxsu3sQUYGIHEV5MJRnedjq9479vupDSII1z0BXSq6Fbwz2CvYxZ9+Jj
LwOzqQ96+ZUJCr/+39OaBPt0A0kkjyLPHe0cvEUFf5i7SziMix8dkISZELu47+XwbH1g2NWFJtsQ
jedG1MMJB/5Y2I2zZgKRjt0wmwVSBvxIUCdh5/zseNV0pbmr8gexX0IfxeVkW6C0dRBMZ0LRTLsj
bI++H5/B38xnYmoMiBIkXliNg50do9MAavwmuR2nsaBkwCUh7lQvUugBZnodpME1xwAwmdMBUcu6
axelzq9HFouimbE9Is4aeTmf+RVecDetAp9C+ggWkMH2vL8ATE9xvbiTHTshxJSEdhK1Tk8KoBlO
Q97TjPPRnlbKZT5CdDypm/ysldLy1990eARrrQTW5ZDz5hG9X8EeDzcf5O2N/oythprTw06A6sv9
ztMcDtqXw3QEVqEMAMWLW5/nyl/qW09DyISbKbEdiR0GQU1LhD9Imo+gSmeFuo/6BJm2dohtzBf3
KdhF8ad/+rFdcBCqH4hgICkUL/haKiWl0amKy3MBibUO2Rbxjw2Apn5WOtNvVxDbRBzmFuLQrHDE
9fSvFolMO4KQ/ozVt9tiUzrVEXln9xCY/E/bTa9rMb418tTI9yIhLKNX75vzjC9++/QO2Dt1vTf3
zIifFmn/oAViodu9arHDsm4f+sqA/AG6GaIQWfcxK+HFhZgy7Dtegwxm6PzGsRXU1aHj+bNdQN/w
Yojx7+sl6hRVE7PIFq9VzsI8Bk8QTnTFrWSQOgv8AZuaTsy/BoxtQpz+lwJJuuwKvCSpljxlZY5b
5mP+asFI5p9Ovp7xSnL4Yhdn3zPKZEDxBdny5ZNo9nA+xPbmzCkkDdm232BBLOD6GMqJ4IAVCSLE
Z1uMFrow79C2ibMImCygDcXpHTxr9Jd9O7gDgXOkBn0toYw832kDq2N6AO523egej2akPoioeHKV
mMs1H8/gn7oMMBAPaVXwIxkuZB3ATSnWVt2VHNXzt/c+MTj6H69/zwvUCZaOocpJDFpFs+jQ0S9M
W5dbHytIcvoq3FaXA4d8LnEdrfsjVhcwGKAmqfQetg2Z/QLOLKufqcHPFCs1pOIwX5DBLCnIa3aW
771HmrxhdzES9k5PkBqrvmEMAzqyZodbKAPPOJnHn/i554cbWkq64cY6fhVE54L87V7Q1qubKgX6
2/uB6uif3Z5TJG9EgOA5Ewj2ZJSkAl5olmYlO14TkcbA1VJ/EmscO3GNMwL/Ge2jjdjKxgQIEWgb
l51b+aggcfrJTb+TbAOPv8W4lXU4xhOfraNYbHmmgzKbKehnLZ+sclhCbuEO6t25qwntK1kk1r8A
+NqLbe+vG+gL2LTdx5MwQ8zCjNPFP1WKlZrWfP///E2dCXzNNcwMntgAN20GkuZi0FDrcHMaCVRV
nXNDvcca52eD8KeSee53gibYpbjtfMMMPneKbCQttXzk8bWDYEh4N5omqMyayYxD+Ev3VCjXrvwk
mhVqKWUqHbPsso09edeMGAuqC3BTFg5mHbsfrikmjpzhXhPH9wjFbUvIFchr8qUlli2wPcfRB025
Htfo4rUe2u5EIc1dC7E4Ru9TBw1mSEUE3sati7BQDoUc8Ian/eO9YmpSZQX7PreOUFWPhAi1HoHY
uaIOZbm0LbvZQRL2sOYHgChUvEIPMikIa0ANzus4aDFGiOSEpIpBthvC0egCvFmEAZSYjvJ1tUGh
YlSH4qbuTn5LgFujOv3IWHe28EX034HK1MnWjkiHehIDiKgcLaFjQKUZ41LhsOKkYEpodmAadoSG
SUHKEZWtTnRiMQruIicywJ5CqD6BgI3K+OH8vWCpGPbwT1w9D1DMntDSHDPTitR2GVxHx+hhuD8t
KwORHVI3Bagaclmd0zNWcNSWJM/KbdtxDqmU07+YUNh0z+/YQNnZejpUY3C6gFMwLWrzo6PXp0w2
CFvCr6pX6EMAOmk76iUwPTbYPllf2WyJdqZFc++V40Tj+RmWtkz/3SPlROllwWameq6OXp/sYknT
UQSoj4PK1FDaLLAL32+lNHRWhjyjn/pQpUol28G1BFMg7igRGlBOqCtlgGlGvht2DjAT3GhLtM+N
cZAPwZNqeU1h6/eD7gag/Fv4ClyF8UNwC44hP1M1+CgtVGaYYuHf04iCFwPGR5z6tXgRj8IIYOIl
O3ff0HkAd0HMTNKqBouisqNVmfAFV79D3wspx5WdjK8Tjoj58DnjGq0OBu35rrQkBtr3t800KK2n
2EmgW9IFNFArYWeoulin5sUoNI8kauoxVz/GJCPE+xcdMf+wQdrHD5JzA9CYMyzIMuuresxY5Wrr
6fWLnTacHZftpULI+rMn3KqafDLzIvfNpfLG+Z+7rVmp86uJBNAiiWrv6VzoOdhVUb2pDZ8azgzJ
HatRwz1Liveu2Yz9BX5BiDh4CgHE0IkDMxwzsGpC2j+z1AEpMX64owg9M0nAW4IhIKT4iq57EWvD
QZkqekA7AHCaqT5/RMeEplLK3OdYPXpkZ9Yi+CQquVYR+LEawuDof8Mg4joPfD99/DE3gZnCm7Bf
q+4PluRSthkbpUaFXPU/NshV6PMNOSTYficxLFQxH3iQx4EeDCfIHq5Oz42NjWPdFRkt03a6GF9C
OtAszRuZeE5+PtcSI92T9RqLLhINqFMwyRwA5RfiNeit6h/r0+7rYvLC18vrEsy/NlkHZzYrjPZD
hqPgDctjdmhT0MN4hP15qMK6jRh+DVjaY9K028WDZ5SMRYF+RFys6l84yd67V4sb987FPc83IMrB
u14faNPycGCxl3aQRajuuVjwGOTVwcyaJjtHdSCR01sW9ouhNtWMFpS0YuiSskrXiSuC7VpzWSVM
PtgRnUhNzEPjHIE8/WFrleuNCc50Z39ce6YWDQCrDhoX8sje9LK+lcZhjfR28sfjhF0afZKWKaCL
VAbMP8CcZnfEjXy+rT1t5R5pkQd/aHS9B3zCqgDvkTASN3aEic7aeNXjKa8t/60BnGkXwBQbuHoX
UY8k6JvYqfvfdjEjjLjvEr5BHoddL/F7eYNfGhO5CRmcmFlQLu2CqTB8W6AvNsa0QEe1fJh/qIFw
aor71zKXu5HryB0TAL4w07pdKoER6+qd7oKyKTo1stobP+AmHud8u0KIauZpZ+2qlmn2pjZCJmjD
jlyXvZepGfxUlZ95dD7aFqbgJzmGaDi6qOFTE3JKykjv/KyixBbmfYLD5p7WZHghcPuDZ37Tx3Ye
dkRegIlWWAfP2iWd/ETH2KfeFORhgArmMaLYjFryeb2rg/WxIXtJpHsTg+2z0Z69CRLwj3CEURc3
Gev/vklpP3g4If+0tU5wETDhuHp2TpF/ZV4jwrHOxfqDMpeGNYtaj5y6mdvEYZ3YSEU8KQoqUMBv
hvy9H7ykbIUJEV8S432P5LbVyPIFzBKxgPviqc9jBs5K9YtOgz/GBXhXkHyi93+zN8PFIQ8GfKXK
ECyRujCBxZ5etiC9x9HcZPT2rBwyWkKN29tOmcPZVMsEFgb1PUhxxxCQ9gPJkhAcrGP6groowZ9J
AzZdWNAcPrxj95yUjt2CRFyaICutez50b6LCXC31bNM0iJZ2od60GY7NQHI0/a2ZfRIpQy3tOem0
kkE9RqSyj3OtiYKLXnb2XKjwXnBBXr1yx5pFhtl+4/Up4AE7FdzwYXoOAr2u1IMG70kTgDThWd6j
zw+heRzgmQjwkusdfFzRlGB05hnMAxEcjfPoDoTh/Mx9iAeCGGzwGMxi5JVrtzxvsLxdSRJqCbWF
8w8nExkLIWdW2qFPltp7qh4Oxz0UgiLLmT8q+MJXI85Fee0qP2CC6lfYuvRPMmed0x8loW2cDRpi
I4jfMPRhAMOXTkAF6CKA5ubHmg9PS6eoZsAFhKEoR37JKfqJH6A0CEE77X5QOuDChNMvhoG25UFJ
tbkzFFHFSFr8YLLVvuY2f4tSiWOPKugbqYL9dde8kro3ZOXiwJKrS4aFG228Qj0b6JxtUJzTQIT9
Xup7yYGNKQgjYZY/m2+FRYca6iNOv3y2cP836PcjYB4kG/B9Ddl6yMx8ubmkpAFU4/syyi3RBjVr
xVlVQNXpGSCT6R/5z5NgU3QcGy19tz2sd/Z1z3sBF2dGknWfnZBqc9jCZ5PmDsN1keAO+VuuXaac
aF+OBQutQijwGnmx1breVP44TkIQvXwOu4RPUEFMNvnQl7ymuFcpk8WnseSmQz7SniTMxc5T30O0
7YkpF0QMZGjcAwi1BtVmT6IJh9ddVoEs3Uqq/ye9srMRe/jVwCyZEc++PRsZimwCglphwz8xbSpF
qqD+eESHssAtVaEAQUw03hDqX4TmRi/yMOKaHbW/f1VxSo8qEdJ2lJdfCALXh2xUXsQ7RKo49hhz
+z6nSr4HDlBhXRSHv9j54HJvdp9skbplOokX/o5ktPZwY+rk4lpFBLdGxlIp+12tW70m8/dBeRpc
ab0007VDZdjh/Vh5Km5I2snT1QA9jkUFOuBDg54BkJRc37P5P/Nt3mM2D9xoPgou+jIMQBHcgzDP
xjsFizD/7Gdgggj0kbnk13kBzrj0F3iFfAiR41PhneA31WdR/NpS3GfUdDU4/MmNZo41xKgRmrh8
vudExixPDJDRlkhao9RRonyaHvW6up+c8oew4gifCarneuRUwl5b8IHyr47i5XQuCpAY/fxvUfpr
sQ6XoZmm13Nsn9Q/+QyZoo3x5OTvLnlADRa9dXFpdL3Dx61V6MNe8g1mxhkj7Od6e6AEtEX2sBJN
pNG0pxjpRVmj3B0n9St/oPNlB/oaHK7eCcEnEJQdtoFusNm+JGNqh7j/Az9rfAW1VB+LG7LvT0k3
uQPaetOjvUiBIMtTmMjnd8fgYp1X9a5EmyTENc5FcMiuRKW4wSAm2OkSEx1ceRihmqrDMafhpLA9
si3EUBMJFWbj6bofg9e1LE/yijAtSGyS8M2HQ+pvJrinSeyFD4/cd14IL0ctTMTJtiyeQD8vrpDh
KJ0bKd/nAKQql22FjF0xV+KxsTQGi3RcxFnKtHd9DLNmfd0E3aaP6kYMkwvFkAShQ42bugoVK4Nn
RFdeOptaBM80hCy4J4bW5o3p3AKlyveMIu/aDpZzJ/SyBC76I876/VWaLp/F03wLMW5e8RUM58aA
H/5ttBCLZLaFJK6nKMvETaZLe9BzZ2f1Qf1FGW4rago0+atAJ6mtU2x+DIm+onINwyYSuBjz6Jnk
eTMx3kR5bWcxkPZbYpa9ODenzKao5XzoBWcsX7Bq9p7TYGy6KvtK7wBfo3+MgL/WN2kcE2FNJ/4Y
vkqtaDJnFrWAhfklyBVeKwL0ZGqadHJctJwwxJpevBkYezamWMYaltjIOns+FlJBE21m+AfbMUdV
TFqEiW7gbCiE66L+9u+LHf/wKGgo9bIWdg6cVuHC8A9bJI93rrexm1TLvbcvTdAYhzqnaPIXhfEG
F1p5cGEf+qnkdT0/q4vBpWRhJwnCV1IE1oKA/+Zitkaraaj/loPTEcgv2Ryomz6qhv/NkmzVBk7y
Y0ep7ZB027IDjCzgzKcvXQLlyYEatRdzrBG5i2OCl+TwFbe1yyMm3CAw/6ndVd4ZjvUJJ25PGSqn
ttyGBAIIW9j4t5sKhAi1k3gAixkmejEsZeqgPaJobjHAeztZkssrXqvWAByME9bTk1HtV8wkDtNw
uUIqgr81EOw45Ig21JZykOEqgFxR+mhybo8ZGyFNtMU4O9zzKkTois1CklXSNf/fSIYvtJIpoiYs
VTPl/2SkLEsz7tDcMZaLXaaFLuxgo3ygyQ7zFI+xQUOr1xybSU+A+xxClDj4jnfZdDUte/Nx1Dbd
aGw0eBLRLyPf3wt6e3U0W5tPE26XiV+CGKRrigsMyp9jr9q1QFVC5pTdYowU3BmFMQf640ABjugZ
O5PwALEZCDF8PPSfBiBQHtDzsI/L3Q7QAP5EYibjzbKQiTsZJggvz4BQstiL5Uiqnh8xtIEytlve
ogDQKzZO8gWbp4/NAQUVReerWe4b7eyy3hepQETFGCNPgjeDZwBWIwg7ELPpTWr4ruVVtBOHmfHI
UPCQRAoAL/4FAdXsRE5iXnaQxPGvP7qwAMxiff6gHTjmiKtVOBERKrvOuwDd7VH/69nGpsoCzG2l
gvAvijDd4O+F0Tueu53f0kihyNLow4ee2zQg4/LnNfCrCBDn6+XhHsk0ZGAErdezgxFFVAMHaQBE
CIwfyTsUfsfO8b6Hfkge+BBGdArLU92tieYKH2Q8tR1biY4QQiugx+h5cl9ygv7jh0V1cCJMAhb2
KO0fXUarO3z9dZ0cgKR6oV/SplmSFRAp7qajCesLco50YxyyQzQrNT45l8yqOmEzidcRUQxjOMkJ
WjD0Yl5KphdM8GwDI8Co4o2M8RGFhEzip1VttFHW6g7mSmVBJrmd9v8vYfPfElL/QNHafLmg1C9t
M9a5hyQz8gKpdPl3wMtKzNJQDeC51yBSmhmyH08M60AwZaLrVvOhkG9MgYlvJ2Z/knSu/31ohmSU
FsCOhU6WXdjqBz6grFpSdw+xsiN/O9W8aAbEjINx0gem180efnUIwvwn9h3TDk+UMuLK2Tk3n/x9
9NQd7gnIQk7MwJEdkKsDMMiLR0HJf4iklM18/Jtcf6z65je4QelKNwZDyizBDWr409JF6OG7h7iZ
fv5JT3gNp+HbhckJfSfK4triVnyS33OVF+Z1h9e28k6t8ya+F8+Ne0KBl6s4z9vzHVv+pvrbdpF9
WSZDdIAdtU5UxR4YfX/A3wC5rMjXLtBZMSO1ShFuc+7bXczn3ji2oTblVqsoidEdcrq7YY6wyM2N
ceQvpoi7Xbu0QHGxnT3LRbAJTEjzDJJHtfxJonY5nV2UXzpfahoMkr+oPB6RnO4KFEzQmRTUyE3z
SQPVJL/hid553EOKj/OmJTppGHdt9/kjvtReqwlmj6sAXe5R6W1uuGkIIDjHs8w5jaY4N0Cmm1n7
0fqxiN1oQEORkdc9N3cXxCEs430VKmNmk6sY3246Mqye9IJyQqpo4KrGBmEvoB4b5uwovOVJew3J
wjmT6n6ZLjEZ6anEr1WvKJ/1ZHJd6v0VLH7PmHDHXQWtVg/jhZmw2o4luze5QZpmvOWYbMKd1Rhf
+siZG7cTLkA0lr4X3PwpOTFYZkq+leUGhwXARKag+/ZxhxT+H9ahkkJ+n2e9/y66/2iVdBpLd100
hktJF0k7ZBXCZ+AyLUOGb6eEN6Nqc0ERly8BJUeStAoRiPEYtah3rQiABNCyhqJehdafgHT/nXpC
DhNGRw1c0ZJ6wX+qA6wKBqpEqpNrnLvUIZ8gWKS0QnDm2PPwFQsDbbFNe1HTzWtdzYGMEtp8ZI6i
xDraAcYcLSOJyFcEDFG/VM5rRvLHqFQtOTkDYAVa7TT0xjGcZGge7y5lQCD2x56fyWV3tIK7Yl1v
KWM5MNQxGRv5olasTzmc6zAeiaheCceTPw6miUtctsIACC28PCmc2lR91+Ox18xzH4EddawMapbt
9Tn3eo7A05YrRd+gGhkQO+jXEBmWEi99AXbj/gkRCJLrO8xcyn5pdPxmsWhtcrsPobZ0Wj7jx4z6
k/OPPHaQ4XuM5eGz77MleeEPVY/LEx2p/07qVR8MMIFTushRpTg2Fddox6Mp+1ALqjMSf03cNGij
Dv4FsqDsE0tghwuZ3l9EQVsidZoxzT98BQx3EvR6Tc3/7aIsYO+nPHwKlTql6bL8Qmo55q6hsfpn
2Vu/tptBh0sxIIXHCJMh4RT7SkV0Fa8m8OYJr2O6RGm8R46GFoNBZ5D7snXKZ8R/5agcVNk4FKQ6
8ayb9k43GYRWyJSTqKU1qw74zzXclj1qP1wwPbyJuA+vQRG1IIVXxbgdN/N2g+mk1WY1gz6tzWs7
oKdidhM8u/Wq+4AzR0r2YNYoB77f2eJnU6PTh27mBKSoD+2v4gfIuePHWdv+MBiQk3iL4c1cYnMh
hA3yhE+9daHzq02nkGQvZLUZCJj2NBKMXvrBt4J4b09MBU7JWOwUKqYhBJD3JzRo87+v/nV9y4ag
HldqwQ0NvXL39dXBTq34Tq6NRIWL7pnfuxxeeCePaIvAxX3SU8fhaaDqrMDTPnErM9COJiKgH4sQ
Q+wCVOe5vZ/zG2aHD1ejy3r5zOClQVwwHtoK0yzwM9fcvtP5th9YR3bb/6HJBmjbC1u9T2Bb0xrv
dDzPrY7vCt10pot3xOETBIEfjRAEBXc6yv7gMTNw41fBKfN1ObvK98iEVfjNgoayN0S06QkMPQBw
LsTyLSSYMpCXnnV4+3vd7Ko4KwLdH4ySk6etP7OynTrKjS+PqP12x0nEM/XpqmPq7bJr1kUXx7tb
ldBpkPySo3kaLI5G47KCG1vgCEEG9+OxN42SRyfXqZE+3AkmqKRb1Va0sUCZxrogChQUIyBEPqq7
GvJ68GKCEiLYMRHtpb8SCHOZs/3yW21dQZe+JQmNB72RNH2kJ/pSk4Q3Hgs5dZ/RIFwqdgRvNeXG
tL8m59LddF8HVRYvyy+FokkCtbPKU1W5S5NJ3dKA1huOHmESAWKNt9OTk1ntQO0z4GLPNIV10L/5
E/qOexRCZmdfO0pE32jMHMoDq3sIjhfAEg91pUKt3jrmh5oJiBA0YfZnLA7bjQw+WCTQi9C8plAH
g6V0EGNmmrgXb+vm2s/ZLV8AAz5JWqjb1uu9BEL/NBTP56upajKytZgznRx6v5+n3y2y04ijvGjm
ikDyJ2xmKfFuBjQ03rR95/Z2eoToQPugrW6PtkYGJzAA5I5e0Doiyc0PXljLOx79kcnwnZvWddOC
9h8r8PwYRcuIUPZLDGs5yHv7DuZp9f7lcAe8mKJeQtH+klrIj0M2mA3mRkogLQmKlxKPgl8Tf3AZ
hQEXANf6TGbdmHRDFDfIdksEOlS3OJKHCgI+QMsdxeMI77YZnBRX/aI73v5IneOLiuYzWmFoYDTy
Juz3dRsMlFe3Frd4iLKdERBRSKEqvNG4pGh0LUfSBX3j89l5cx74QyCwDFRXre7kawq2O7fOKUZ3
wfVAOza+yWRBhnvi+M2yHYZvWI9QPb9rviw8cMO63yY7He0cngWKk6uB1KeiDxv+m5h8DLYSzvhl
zl1e7Ps/Pmzn+SJ42rnE79h5r6zbn63rc7sdc5vv97LL22cDRy4vLF+fPvrOhHuWZ+Rng61q7XQk
nRXaGGOBuSOdcdajldQrMSqT85/hlU/ueCEc/j+PTKTDlLmOOEJiir5pZS+u1eT1M9Qz0L6c8/2b
fxoz4XkxFGbSYUmccCA4ex99Cm+FAQ5uVeHkbin7NFlf4sjKc6ATI7smVFdAU++wPedcnve+CeX0
0NY7MC8pUBNlVZZnQSVA3C7eJciSbYarpxZXjZ9Si9sHNCGIL9Z9gF9n/9EXPiFnfchBzgX+lABq
70St09MS31yx2Qsu1PuT+hNo0h84mSjIGfAMclEh8WXgOflyQe6IIPNmT9tc3dZFZp6S0KHhsYDs
cupAt0VqSqgJINdSPuvxgNN4NixIjUGiWHlUfWIXJ2QtyCIp4AybkdJieSy9DkTgnb3RrqZbPqt2
imgUEq9bzrPOU4AE2Up3x/ib0sRO2qa/198gpFHIAfbZqEnkfZXjM4x9yyNO957nhTdapWANqikT
JrX8k1h2LHBBd0P5S+904TxoOrUhuVJ4Vj7clK9cFYw0O7/7xl4uh7mRx2wlsIrMEHgC6L7aphu+
jC6/EoRkCsvvhxfzNxFMZihX3Ue2AyP76guPzznGb6bSYO1nRR/HpITQLzPznALF0DYtlu0zByvu
nY/5b7iyPBy4U80ri9FwL3rqx+AHGgsL1cGFxIR8qpdFaUH4ivXvSIwdr1z/FUo7Y2sbfLWZJi06
cnYo2UtWAXnapQNV2wUeDraTR+VtNwKlH8btahEVzoSaFRFwGvH5rtpG6MKu0G87eD0D3Vo1P6ts
U4WsXUy7TdVvrJi9Vk6An0t/9a2O4Vu/TZ57G3MLVg5ZiEiv30ZiNpr0cy5+dvblp0GqmX6cRjoD
5YPaNJOgvN+5DMMgQimoDorvGoQzLw8+3LjRlmGHRM56atprcCsf41xZDmTCgFwhb2tGWMTn+3Qq
fiZWJytWZFgP+StdR0nRCYOw2gSL0MlxFVEKdHnlBizfa+q9V86krxXtt2avS+8wy5bwWj+IHMab
x1aRE6BDAKK3soBvkGxkM4lmcskYH3B6qNzLmTg2oCT43wf4las4F7iFrvTWJsG+qjXKauZBDHMD
w7ccEegyAx1Jc04DAZHVsmfy09IIMVmLNgtih37RYGMdh8DgnplwXYf+0b9urowBuAYWkIU189Nm
7jXgwTnvQNVU87hhcb3UkQ8xjbfC5lQVFqFFBG4SQzkwacttR0v1naVeP1k44kio6704rxkkaniO
cE2NBqz3KNSXRPUHdyQNnJOka8D+ZgtN7FybTZBmojchQSrkaU1HtV6JYVwSbcXB2E/7VxPqamlC
4/3xoleeeKZX0eMmHdKBqgAT2kiNQJYjpSBx0TntG9aIMKUqpwYp0et9fSFVkaFnL5SSVxcOGRDo
UTwX5LswW3umVarZS3bcODczM+y53JYDn/47HEAsIEKCtBs+ZVC5PhICPDmkJPXbeeuDWtdqzGEd
AG81XsDlhzeoaUYH/OiGXRe4asumgYdN7jsO7Up3CYbnoBOBvp8Zmcpa4UpxR+gMwyer+xH+FOkq
BX9+0Y0plEpXsYRYYedoKx+emqwrLrE5Bdy4ygY0l8/0bNv9t/ofLUzmitzXr0ZOL0ngyGYSjOOx
ijTzdzf5FUYqxBdT65gbcMhlb7Q/1raanKhRiYsvaPu6mNYVSp8cYATMOqw2cd1b3YK3UuyTX/y2
tGyCgZ95dLkMlty3ZIzNNpA2aVaZcV+WSQY2wCjjHvRvJSy52kyYu6dy9pj280vfdcaFqsJF33rp
f+hD2isBoxQkzSH9ez1TV3y1uNLKg7ARFKL7xAB7RxhApZM4ne5IjzIG2+reQUr9ArAsjY1krLt+
yWKrPS2D0M5vGlrfFRNJfWKwCyWC+/eVKzg72Cl+M/jejPWX8ShG2jTVHVv7K9mj28BFsTQwgsIJ
hHYiHQJ7HWik1NGhRLXG4daRx4AeN7GZ/DDQldudW+s2YbMKONwwlyQfS3GExEK0F09HKizrj8BN
/5TcW33Oy3kfcnYdmyFLq6Hpvyy0pGsHTwga0r0vZ55BijwA+e6jsVPEESNfqoc57Dtbg0LrrCtt
GM/I+Bj5dHCOCtAYP9KLAQBGXWeHp7T6fcCCkL3mSv32GkWzEqadFmRi4z9DknrS7wS49iYe7BUE
3I27VX+ifOWSJzU+aTc3fROLFQWatSSfD5O78bg63r8JcwhI9jJscmlrb2uGNQvDe/NnxCTR8sUR
IBW9xr87UDccv2U45Mo8vNpXMP5BaE0b8Jcz2tgzyugox4dlMuidKI1/T/D+bbve73+AyEttIDK6
jFa1Nn0nPWDZWYkiAmPlHXW7Bx0/WPETj3ufTwDD2PRQyalPLegm1IalkrmGFZSMigrHytgvWAsG
0vKuc6AIMF2JHTO67mDf28jxdHXJEVf7vNID0WcftigaRyBr9P9Xt+VMavVUW3y6MF0XP5vLrzIT
o06QkA8jT86BLTMceZhGoP+yhGSgAiNfAVNCuus0AlU/3W4538zY4NPThgAIPfgjaujwOOpgyPH5
xGyb8sb6t2hMtN2jDLzQJ7fvigfzQ43G/WEsogSP9aOEFR2I5RjA1uM9s+nvfvvX9r+Ujn3LVnEi
lkoVh/SVdn0s0ePC9d3VB4Hl2CLj6L1mwF0TPi8hmiG7oFA7CN/y6+LCbxiDS/2VSb9DHFLtz0ZS
IjtYiKMOnd5/Ope/OcOXzwCL0xE0KqoNkIvqjNzDJ4SW/U5BxOpqIFYRnsdBKRf6kiqUbqkj5V0i
rj7xo3rJvdjeHJ/Z2gPqNdwXO2kkIiagUnszsetfcDnmK+8h8QACuR9A+kQPInBh9TqxtM6pTQfR
GqJyHEnt2MbQ3sA7nCqeq1mKqF5yh7FEcjyCbkDXIv5cBntgzzQ2xnXekh0uJJ9jch6/97qfWBIE
IE5CFSt/I4t4quXEc+lZ4Goh4spFigIUAU2SyU7MfAmYSh0bQXuaiXguDnhGsH+6O0CVYOZ9yA2N
Ky0mjbm7iM0Qmsx7Ik4kQMHcVDLZCyr6gD+lMCaAYeOn4O8qOSdQxQdscplIm4BSg+HC04IZBB9n
rumybKgFbjnYpfmW3rpnqk7x7hpP9O4ztRsaKN2JEpuO7CoaqxRI8u3z5570yrDIJniwaXmT6lGl
wzK3qcxRY9vA8eT4CaeayTN8NZcRNahOMkgw/AVZ34Py/Wgc/BVTIHmk7Ih+vsitKkwVMNywe3y4
p3hsxMGYQzy4TycDn/WbpRGbdD8uADT/j83hEAZARC8bVCmDb2D94fc3xTqfCvVyOeTGqPZ/9QtF
PE+vxInidK7BOFQMwvTcKVgyC2IXnOwqjw60aO9lG1mGf8We+nVXVY6KQVHl0G8Ur7NPFUEqbmvq
zkpurRWraLIni83CsHWGk/jygHV+vkLK1eQdaFdJ1aj0nVeHlFbZwV3gTYSnEbwTei5P3aJfd8yL
gUygJbrQkmg5BJ56kLD4ydE+ywLnIHwfIvNeMxvGxun9CUO+TIoXSqT9xuDEhVTBXAQjhsm6u/n8
IKhmxTuxYPM+8s6VwA6boB5xBbWf+wOrbOoFRux+eiYbUxHsKHZbbIq5gY3m2/YG/Q8ZyPUeQIfW
ntck8ahOiFgDXC7RNeX4geUduwcAEImYHLibNvTPxlXr9VLL8qX9+JpxYoiTEKECUMMnrukw1WfD
yBEgpZhXI15vNk93lg9XtPWGntdWhrgHot0FW4CX3mSCMGx/4a6tvoAGX0d8DUiHupTDnCZsuRoJ
BYRUvlMJkTYIs9XbBOxIXgoYii4+Anrc5pHAx9iFKqsNkCpDD/8hgoPKCVKEaFk/Cuc9O0otdq93
RjDIP44h3t+Cg6CPHS4FunpYgaRfFTWXOu73gO73cDBZujTz5NjJe17Rzi7vWoF52v27FTMWGGeS
IlrPpF1eJ1pOAhs3zc+sencjtmuO/tIByvxRm+U2KD/RNSb2YQTjBtSw0tQxO9HpQ4xf8BIIlpFJ
BSxojry2OaMkLfsPNWWHfKXqlIuZPrIQ5E1YpSwf3+kvPCT49R5bgskpoJ1yRu9rf+KEY2c/TziO
VzKOPdvM0GgaCLsEy1Z759r8EPqSe3Jl4HRJAHKTmh3F+tmeR+PRj6QfpTW3zNnxFhVyM+Cq7mH0
+txPcbbr9QATOtSianLghy3D+2ji7jdpxJmaP0rYyQoaEkmJbuEOqjqQb9K8V0M0xKx4nZzcqowd
KlXMrCZd8OlAly3KhfJouK6AHBV26+JkIZXXy/jPhBrgKsgy3e75mjs1DjZyrX1Qz3bcVT6ajQIc
je34TMtRcMbdXHuZD4jaWa0ThimGxONKL1/PhAw6kvGDZg8WIcOCpIPw+vlmRM97dJotEWQdWMhf
npFKVGPyiczTnNXlI7V+VbEx/hxjV7DKBgy3F4uQdpu6ZYIWcG8iljohrhIRMJFFpvT23hYuAeHh
HbXcDPsV1rWPRCqLKZ3iTUAA7lmAivaCwv87g9AaGoNX881LAoNBkbLggtFBnYcpdgq+vxG9Kr+g
GbbfcDVo+0FT/vrh17pNzf7Rx/MI921Q1JoSyL6lWv8OsNsSxb2y5rC4V7PdQCYhHdTJEqDeXAdf
oRsYsyPYucCJVWwAT2hfNPqvpJ9S6CyrIeIFxsM2MFSoYHnx2+2rB23r6g74gBmF+Xs63Hyd2wZB
mHkg94Iujvesn7cEyEwFqYDH5ZyGnjSYeknajUpAMF8hTE9Q0q4VKl+jteSEA3pged7WOlH8C0vu
+JMcya1D/ARyoBcQkZfCvYKL2851d+ahzTQhYRbZbLRrARwMuwpkZ25MpNx/i8Ir8n3+fsH6aexn
dCCTB0XQfqNRlgZ59+dhngKhAs8TbE8TGER4d5b0ZBesJc+RT15NmUlsbOufNuELxM1VV22R7Qtx
9gokeTM2Yj+a8JXMZPqvPc/bm7gkjQFYvteCwl9iOku14p8AeWRNkOn/KO61RLaWKYz+4N9sNRyd
PlSk+jotSldup7N4d30x3BPbp4u3j6aS2ZhU8GBepIuHlaIfk8ZDARWh3ekswDZUNqAIsLtyWn6Y
HxK4xbfrxtqdpv5yduaSdf7Ii9mGD5a1QRxyOx21XmDRTPUADrtgf45dzkW2SKYbtIXGvatdCUgY
4KuA9kZnnGn3amLaXPzMZxtzrScEee8PTFw8vLSGXyuy0TM5g1Dy8Jb0Yj7KlN9g4Lh2uwPSBuT5
CLJ/QXjjcoqFXNVK1o7W7YQHvVcFuUk3cdpwxb6iR+Yw7isOyYJSoBPzughjBMfLp7bLZZ11urif
QZXO3pgvLibUvh1UdmZsJkKbHaiW+xzE6aMf17+QhgYlFY9hDl7db/MgAE19Yk46WcCLzBDaknua
U189D9hIVNwUVIws6TzJdqwZ4MWHc/7wYoQwdxlGTqdYHwS3tTnzuHRiA6yHeTowhJtQydM+UR88
AvlO2nrQVIjKAeVHZ6bq36UX2FSVnaIGNtvVB3jeQX6+LLSftaadqZFH4583+Gi13k1JfvQiyfz/
HqRe4vaRiFR3e3cSSxqs8SfCvR8gfoy4syU/0xOXxIef+c02FJv41dm/9tAcO0B4igkfGsr0Wn8H
FUx3iI5wasn/D9Gy6YKT+Y6MERDdbUAPBannavNCRtrbg9+qUbFIoaTaGD7weGC5FcxVwMBWVmGS
tzZihdXZSuQsJ6eIvVpiBagrrHpPS6F7e+ACGwfsy7NeaGO1HfM0IzgFV0eMTZ/dWTprwFndY56l
a0Aoz2539Xn0f3muCtl+CqOFGH86ZSUN6E1MGn1fj65e2EoKSd9GMe+h7Js+g+xwMjTklt0KH4Xz
o+0giwjvhm6R7a/6CAb2v3aX6Ce8RuuYMwRLHrw/5XdMwvyhhnlL1d3jKSM3fC88bMlp+Lyz0VXz
/fvgHiwnNfydrMDQlpFGHeqnbIa18R/tNCqnnf+yY3rKvmiRkpSzhhenT2kECQp+qjVeSZPpH+5X
i6cSjBTvMU1YfsGzRSvLc+KW3uaJbGJRZiF3TcHb0yT2onVItbkskSWWiST+YFPmm7AghKnVLt1Q
gO0WdYSj/526qBNrSwyKu++zxDIr+4Wi7CSpCQ5C4wSy6zikbshGPkmkAyDPV0hM2a+ct0N7FImO
P8PR0E8mp9LR4kHaSJMhoFcaSnzXPWzg7jWSaLgkJCZ7h5W253Jb1DwcDvSAnS4hVYT5S6DREnzg
dyVvgMBBYkdGrCMzZMkv6FbHxppnNpqNRKqm1D0qSsEShwkyh+ZGpVLv/edG2xVcB3MZx3sMzbJr
eqYoB3JQyTJDs3u5Y5xHu9qAd3irYpdRQz5zCFumLO+J7NhTWaLb8o7KGluXwycN2Q4XmvbatGpt
hvTIbHkhSPnnBCzsqyDjJFQK3OF6aG4PHU2pf3BFxGvpYvzl1bnH2oFI14J2msi60GLOWJnw81Bx
PeNwx6cHGNjfdhPElb0+LSWIUkiSnJV3LSVdPHc75ZlSTux6Q0HottwhUhRRu8hNkLxFY+BK8VQg
9WI+YwYsHz4qawDYZbrOcgC1HTmK6JN7Eo8gy6yyI8jlaGOr0kongd3Jr1KBCgJZymhzftmIaz4O
0Tll6xtdoWOfbZPk1x2k+oBjLayCaFNjvaXBDvvwE1wwH7bL+EUt4viZZbC6BICointqNhaTq5cV
Gp/1PEFGTfLj10FQZ/cwxIn/w76JIDGIcVhKXNvAhH/YEsTQ5up9YINKqNVcolYGgTDkCzY3P5Qg
aoeyJ3c5ybHQ9FZlkcqbEQck9dUl+hVc/xr7gLDNG6Jae9p9WaulPHblnXygWQe7Nx3/pcHbSq8q
Jr23dr2Tec0KDvy55PWlr+nTGpyL7zWXztG07iI8rilSr130ZtseK2yjkLHe3a9F8Ns5rR+kZF0E
gJhShYxdUeVnofi8TG8hSds29+DE6G4QbPJP2KX6PkRTLgAT4NKEDyb77pPQLHCDsQJKPKEsM58i
G5Y46Tx8MUASB2RrsznpbWzs3plz5x+q/+zTkX5bz9n8wGd9fY6WGYow4VdKD2GbJCfnQ5Vp90PV
vtT8daihxwMo334aA7w6KQRzkvDd06uHWglTPHZtg768MWfQM2hXOKgYVqwzhJk/yLt7JLt+0P8v
qL2ZdMtB6QwFFBFCOMhuHDO34J5ztzxeh+JvstWJOsIM7Xk1MD2bElS1dyDvNGe650Z8jc7ghSWJ
is3bjiyo8sJuUxA8CsicooHlg1BiDBIiIKKDpm0+qWJGYsrKcGtX/kUkO6vYZB7/kr1hrBV0Yosy
zuTcIfj19zfJit/l78dHZTQA4etPluj3hLnMKWBvolhr7YBy8YY20xpS71ceMgz6hHYD1ShWO+ux
5tJ53TZvh4lKlZgIhA9E4EWcV9CnnBqMZJtnBFiDswUNOVvs9F1IN8s38ssHeSy8WPS2UCpk6WFN
JdClkJbIYvntYzC6EEzDLenUFiVNS+4QUvfErdJj1rKSHUJP3cimvMXbKQyEdM48l7JjoDo6dWRz
eoyzG7G2Ba4YjMGVEvoYIWpxBqsJjmC+GBlGbpi/OHwpBjFj3UsbvZeKVUCLkwgzyDLHJPGMS3l+
ME6LuuiyoM0FPDe7E47bAB5x6n7tS7vNj4DIao4MuwDC0MYIMdR8XHc9Ivv/YiFHysevEZ6uGJeH
dTQt0Ukkdnxq7dayfpSluyDg5Z6USUG8kHf8TOig825NHAocAD5FQ7Myo5yGY3p4bmsivFYTFY76
y4QXDLurbOsSYZ3xyfoXFUK2fE9+qutN+8czlhXR/v0Gtz2EC3085JcyH8yreUvpL066iMl5e3QI
s/obfTncDFL/z43udTcSV4mga82Otiy76q2p3HlEGdkhRYBq0BZEXxGf0nBNTYcn+bu2RV3mkld2
LcsfShi7D9yzDEAGIt7zX9c4vwLUikAaQT0aVEa8/fnAd962jOB3/DAkBVSYy/pPNYMjmUyuToP0
hLpivvKO6rr4PS0mjTqNHIPosQPNbrUFSkANtqGMsgEHaGhtdDdvWBA3iImZ1bvDO5vOmYG3+/K4
UGrWllhn+zDnoTvODrdOdjBzsImWLA49evMrYYR8lF7FNZSe0Nl+NMzmkonvpe3YpISv1ehXC8fo
jKOOf5q9v7UiIbcmGArFxeGsxk65z8cqEu7RjzCXG6C23jUeCPd36PR2jEO0U5sjrqZXUXMfxYnN
NU0gFpsoO+bvhI9U71H0s10nIoM+qHrCnEryXgN4UqhGReOStNtAwPWIlce1O0QhU7V2wznvNUy8
orFziBsHyOChyxCJ/+EuJRpjoM3cT6FqAkcW9XerHDFmSIxkmtCW80AP7f1pFAdGE1IVdE+IgjXH
hPq3QvRQ1pxBkMeA48Mk58dmwUoIPILNcW31R5qqwoiiqL1NDEJ+VvpLqVV3V8RIDCeeGBL1dXnt
+4cm5Nymqw+kVoGR928ZEYySkzaOqXy8owcvFZWYznwbUxHrw+gQxZeqa7yiAhsJTJN9e5Cs/qW5
YeAFYQIPmnY8JgpIRMu/d6ncAsJ03EKK4bhrPcysklUWMnPWGX2ESDcI12uPuBVUmReqL2AgoB0u
UIPrJ7jmfK3M3OfZt+o9fVpGQNbTxUcbwPXTVlgTiO+eKhQSMCijPFbqJ02Xe7rOuRLJZfrpJoPo
1bUa89EVUSUG8OkqDGj8dfJR9cxzDLMsYa+WvSXKcaW70Sxq7UR2NVVS48UsMsXhYpHsn5y2O7wX
q3ZxkLZ9ii3WZ8MbHTcdlW97/mnJswAIQ+uJAPmo66cHoEoGL0DxE5hdNIADjz8S4w4YuF0s91ie
YkBMk94xLI53THr3a9/Dj/TuayBye4/SkYBOYnYli/0f8wvmENI8x7JNR6gnlML2ghaEZc3TmA3n
VshYgEjyvqwm6fS7NUTtRggHrvCGBwgl5SsYRI/DNsbAN3ntqaytgiSGvCSSdzI4LQRzLj5DiqHE
fYrBZWwoNl7radfEFszT6FgtYR3T0+JccNinUhHGLDqQdOu1nYTujoC/NzFADivSmzEqCi5SYWCv
fqK4nlDo9/adhxdTbTOad1ZUACdGT3R6zU/C+xBmsefDU2riVP1FEkqGclkZ3d35H7kgGKyNHoiH
o7OTnRgA6Weu+31sLxdHFoc4NohA2rfP7Dkc3urZ7NBpiLdwpOx0ZeexBEaJrHHLgqwFg1NRV6+R
3yBJ4KBVjrZbW8EDw12Aw3H+KzTNSfccSUzuln6mVe+PCKfcEfAHTgrMljKD/MoaBeCI+g/xKarH
f6R3+osQyCNoS/B1+n8B6BacPbKlB3CK1xHGHBsI6f587lpLbZpTXeiKl1ztTKkF4pYraCHSISQp
E8fEzRKOA5ObKf3EqJtU23KD2coayQRshsb8hhiBt8bGg+3IAerWDZh9O9v6hnOy1t7qrG81lpwp
cHaZJPYV9zj4/CsJoWwfpq8XKBPA9ZdxA4F4mTdUjte7rxWcqC3RWvcigkhvu5W/7DMnZX9Sjdid
lYjLyTIlyT20b3UMtyAybTZ3TjJoEV5xN8b/lUDjytr67//IOTUeLFvRfqCpZWjV/hAS8JJDIGD7
dzH5mUSo7eKtixqp8LeSglXScXgQwD859reB5fRoHhiH3f6nsf63//mlIZwfaQVUq7yIUb5fl5li
tr4JVPAD3THw7qVCImctTZlFm0qnaz3dFKVTRkkqFiH7FFQPA2MNRXQ/1LusQIxYcve3Rp0ipO0S
4ZlZayEkVq1mkAtHoTbsnWThn4eCAgJofk/mGMxz0awsQG5ABbsu9En9lo+Z/eEJ4pyLkq5SP1o7
06jgEEv2MCQHxiF1ox5uO9ZlU1sdH7ZJvUWM5NwrJneVKVPznCerKsaydZFqGnA4m9eb2H1luZHh
P8L3504pL7Nba1uffu/QY6/7r8e9sHoVWNDoDjvHMjYMm5VJWWE3PTxay71rh6RFrN8dQocI8aW6
gReZwWSjKLatK1AiSZN1pU4AQbtubo2yyTo3rAXDF+R4PaiuuQ5OcsufkEBS5K5Xfn5OIQkDNM3v
IYFQINYB+OiKFPkpQdhmr3e9JSo6PUfLH1f932OGxCNEtHStXP/9RxMFDADxa1QDLla6EPFlMPN7
2AUUrGFLx8P3p7Sq4D7tuRt91uw3++ky4u1WR4GiceibVeEaSov49VrbQc4O5YzVMZ4AbQEA0vKv
cRH6n/ZfXbfmMUm6xQ9PzGRUNaPva1pVf5C8xUoTxuuRdNS9/wwjwkbS6kkXDvrgiYXystpktuZj
NvpFtKsm8dg/oLN5TFaDOcj+bnch8ZNZf965bjyKXj74sMKm2rIQANRzgESqc4wX8SDTDTgn9LO4
w24G00neTYQBw2siVUwH03NpwSuy47ShRDwM8ZKOW8uJIhtT1CgTwVsC/hNVu7ofkonNmSXP8J8E
rgPo/+LSK3LsOxH9UuIphjAxXpUSM0+ukqN2rsHOd7a/1xuCw4o60uqswU/QjSz0ITh9SPpLvCiK
7I0FxBEXBUrC34oggjTdNnfXzqSEDbvb0CQe9hdhlXtpkL9arqQ5kj6YRnY6Q5WrI0JqgDpJu5sd
HfEL5jvAdMCvuV1GY7ENhBTHEaZgbS4QlEeb5GwEsLKJStPsotxEEXBjSxYfGut2swLaXzQzf+tl
h3rNpnT/RDO8SsFApvrt0qwUlup4eCRFEGI8ye4G0PWlTG1Hl4zCwqRdTmFct7QXbtVb3aYRXwDj
bPix6hBQsqnojozri5Y6+CgaEmOnjMxsvIkuifSYc8TRHtSi9cYfVUfLNm8sKqtrNeGwTv28wBuK
DDCcnGj2xGukWZberk/Nb4/6/h9dMI2GgbjxPfJP3wTiHT9OgSuv85LP/9YT4b4qaEN+GFTFC5tY
7TdVjYzmyKimPV6iLKoqkgkFiqyewjpS1XHl2eXte7DdqzsaAkzGkJARU1yeBStjfpKVab9jb4XE
KtJPGCU3INQxvl43oio12kM3FdAbjdXEEXG11Gk1XnnIC2/LKX+FitetykGTV13R7KM20fE7UETo
29p3yLtOEQwTHpuRZHRV75nA52++rGk5iodWdqr30BnTsQdGiTQZcW0T/7VkRH8NviL/XlJC1nuv
Wjw36QXbAPMna1JlUJWtwnsjyzJbUO87SgsryD51QwyyOGXdug4gtAhqYXqrPQDRDm8Kr7kO/MY+
nMZ0P+4Rs9gmWRWzIHjwyinm9QUv0JNa6qBhuvKdBCpcSEOgHYln0dWY5rvseJBpp4KgdZy8O3EV
JDQs0XT0rJJ61J6DxGfMhmrCU61gpOfCAMVkH0oem79Es4lB6ejHZ/WKgnEszGZ/BwNsCAxKYLgZ
jbYQGk3IZKWHpUDbBw/HYVDSBhum41shHQ47lvTmBI9NYZ9QjuGXgal0Am7+kpPZKvhrg9/0xGdf
04PKCuz9m2G1etG01hrG49AXIyJYzSP29JuqX1L8tYDU9hfrsGEOrAWtR1iu1mJo2VVm+43nDiQZ
ZdLFJOReSkCQiSBo4cMwi8kLaFOfXP8T3sp1X/3VzDkJgSyhTpyqYCgQ5aHMpX1EX/lrWgPS3VHx
CX8SbWKGcnPFFQpy0TXL9UYzCQwSoOzaneNlteOulOBonS5r//3ypGdcVl0zCDK6RZtUPWag1Y43
/6064kQsm3NBnRRZHlXS38KjLlPUbRFZU9eE8geocL9aMzpFS+Gr6RQ37Vxf3HbSzzt7UjMxeA6L
rnlEQt7PfeGAAmd3opE6qeeQCAs7L2ZRxc8ZBVXZ53WNJNqBVtOSZHOVy/U4ANdRs4ON96jurVvp
qe8F++T612Sd02R39UwbWO7hQZVaL0pR8M+CYGpkFv6EMHdN/gEqQYZ5EC/uQOsXv1+jpbBE7UDC
d1xkF5YDtA/HwP3dfaIXxqDoWDUSwQnCpBAUvNiASHDFSg6EkmK+BGb4De+qyvPl8xqrRATfb7oo
3TNav+1liXRZCSXGVvF5gy4XmIzxgs91F0+sfQWzWKtzSIkCctzg/B69+/Cv7eIKG/eOQ0SoajMq
/Lx/yNXnipH3Hh5bxTrFWmrie7DCo2rbx8vx3xeD6gsAiRyncAPRw4vSluzsMIsmNo2LNalFmQNV
IHc80wLy3jX2TbAhswOenEZOe/L9eqX0clVVUxpBgguOXrARR+T9z+SX4nIL7qW5de0wIuvikSfX
+m/FRyHmrO4JlNRMyGcJH5YuVCHt3YBAGf1PUTvOwnjIf3KtkjKyRA8e+y3bCiRDepZAc6y+LH+v
cbRstVYsNpeIx6FumYSaAwlP/sBQc1JAaMoMG2RW/L0u/a+IR+skAs8glBnvJ0/IVinrfe9pWzSn
YKBwXmp6RsnCHYMSYKpdH1ErnFQMaFyF55PH3ijmsP15gPG3V16PvCHibuY3Gx9HjqRPpqMh2rQc
r1JteA6SHdYpyI34eyfPhZIL0GW/N2aDZnnwGjkPiqddXnuyP5SViNGkkSjqdkxrD4C6NC3CUgdL
6hovWVkglYZYlf6oLrdl2ied7yZzMnAWe7HKdvsm2HvahBd9qBUUj8s5qlzDmjfnT0SlSTJv1Wkr
IiH3Fb6avF/fZjcs4WVkbOPomufi9AjdNOFe3/x3UVC69Rp7qEEw5n+f2vltaX5O2RSuFfv0t5Ra
a4x96zLHclUGCA+XG/p6CY2f77l1Davi9XT0IfB3JXTpxWJz3azL1tzfZdeHfMRmyh5MS2KGOPJk
qq7HcHGJx0fubC6fHxIQFamRJuG2F5lDJgfAVFsevI3JIX6YDbjp+rUoVvwddTOmK77f4P6PGY70
qKIWM4410oWZirE/t1SXzOCiQFXy6VRM8+mZpKE6ekumeJnxfn54E6hagc/q3diNNAnbD+fBMK22
YvdyKueKrm02D+A7x11bTu6iFxQFY7llZvc3XnFNksM25onmnlIlBhYMK3VWUlhoBWhOuGvF5NHt
m8eMMGrLC0BC6rdQU5jsq7xmclD1W2FTQTXGCZpFzHZWQoBiz/uun6PF4rtbaUI8jMbQkDrdTgzA
GMCT97sxh1mD/UY1FCtkWiNsycXHGNDCcPQF6lQXBSoIuMeZTKQF8CqESWW1Blh/Sq6YgagPxqZy
aG8WwmsLpXau/OWjd+lEldNLIIYkp2d3677cQsRKpnWO9jf7UwBGfMCTL+0C9GvzwS1ZHiNH4bV3
bCvqFcT6tLiqVGQDNBoO+7nch9nLUYz1GgEQAJvy5zlDK4BnXQlPulEXKrH0PnWMU6BDvOrVvrkT
r5IxTofX/e6gp9sVUOf9rvQaE/NP7rTcXetQCP8FGIzikDan7tURbOY4NQ701AtCx1/8RAkMGmM5
r29KnyAKhnJdVmvsm+abADAsXJdr6iX1/mVFBb6PKSzTLqo3/YFHFTTaZQ10BQtpSGNBC2uniLB0
vNSpTDWA1pAsnatB0FJ5eyKbUSWaHTplfBbikzLBedg6GoQN3vEmBgvEdsbE40uXyiQ5PaqgDe9F
QsupF8Wwpai359Csgh0c1OVnlgq4+A3mLFfT2OtrfigOvNxnjIcu5waX7HvOEWJr2Jp+8TEJl4/m
S3E8hKZCLIXPWiMGCm7qenAL8WEoP/MZ9B9+1t+B+X3d7WDUXusU2CsKL6pVWU7OvmLAtgxjdLqN
TprNKuxpFZnRuIebNi4jDWNTL5wDpm4cKBTP0cYe4upgfJpvz+mI17sUtYR7/isw8QEOD7DKmgTt
3qnG85k94BKDSl4bXzVaTShcXNbALLZttVtVpCW4XJy3eSR7h8aONHec0iqELrDKHSkSUaJHQrWC
v5v89Y1hujHrO0+SxnLyVl7N9d4un3iHmbi89GDr7V3oQNZOghMyPU5BtT4Sl/XQFk2Y+B5IT/Ow
N/PdxRPv7HL756m+6HWUs+MxT/HpEM3yEaHfzOtMsPcdyT8I/f4FnBztX3ECBMGDvF4YrnqMk6sX
DO2lr/g2jrb3BAW77+YaqTAPJf0pwgUfP8ZO0xDgpux94SEc1BR57/gqhrYGFy47adZfyXKlywcM
P+YXKrjnvJHjoUlDGQ9D7mDBPoCJQ34X2zq0Zwrzuq44pv7EL7QHd93ijl2EgZoJY3AuKBs6i8jA
ka6gUdcVgU9JJGpm0k+2lEBLWtWPGURx7zyrRK98V33OZRjPYf+zfg7m6qxrxgwtGthmuVMlinwK
dVsTiCRPPL6NFB2u3Dykfh4o5Li8D7RsUGiz2IQ7Eq6zNpZofkdMRXA0aOpqu7ItnA9bo16teIuS
zCH+N0s3DikB8fGn54truza8yfe0+wiAuywnS6m8C9sPjhqyJ/i9jszpGys50amOIuYBwDUxrxmr
5IwNU8ktvzhcydHn6vP/sTVwua52udysIIiWbDMovvMVFnGmlYanFYKMMoc8W/8fgSDyQpWORCTG
cV1Px4xvAmU6ghZiQit9YB+PwnRCJamTtYN3etmgFWA0TX6H8K83IDgdlh72zNHng8YATUrghrMh
uLmaSrinR49FAutkI+3AjmL5X92OKvdCIdpc3v1eL9B2ewseu253616jGbiq0p3Zg05o8//g0qVs
CuuGchWQw9GBAQLkzXtgyJ2nZu3zP5d++Kr2yYjlJ/gyOy11kpCcxG0kIGz58n49Ed4iZxxR4p+N
BZG0T55cb1Ovcohv8iUpZqgscr/ruGY4x27KQRawqJbO2UP9j7C85TEx4TIQwv+r/+q4kNRBaCV9
U+wq87dH4nJ2lszJe57RSAtVtdOjXQH3fVne4+sf2/W4T/U/KJORyfzg0phWzYO6p2ndbL/Rr0CA
l+pF9YVJWjxeejek16sNXDXTVQGT6vZOvHU5UR5pQwrVzoPpvz2/Vw1rHzJnHf0ll2dCgitNwT58
GfgisX2rwLzEmFz0EuChe4Q/Auej52Kp2+kZL6f+huwCn3MR7mD2i6+u53/FICHirm/8LrzkEyop
FjCKMGmXWMoerjjn5sDYjVToWMozu1OEXarMBoagjhTUgRPgG48GWr81qW5rUXwYI/gfPpe31w0M
Ds+kviwVhCuVBSK7+nEXwLF+SsuccGFRtpdjsbbVN8I3iLrjkE013YSeEZ4gnFNiEi7hSTNbnG5t
f+PfRwYo+NutxdLNQQjGzXhVk4AS2K+kwPFEpekIA7F/lVZnH/ugLL2u9qQPV2NUMckBlXa6YqOA
SUrMjSaPDdSUH/LlTwMJ0kf7COxZQFEUBqYqSg+rK+eRLNR82exUgqm0Hgs6vIA8aL/IztKRHkyk
twAZeSqOUIOqSlrfjodNnWjkwvCBCff3Q7KXJiUrRbpxpBEgj1zgsE923xbommE/bFnY71Lj7/pM
/Ue11rucZ5zqDIsQvpPAunLa8tXb2wBzGLk0hxcrdw7HcU4bzNP1xMLoyiAS7AlhJs7zr8coaabW
0qumNco32y9RzmyH5dTMWVAtdbRQ73RjNj1CGZv7tsuzouTYMgwKhqR7/DWWFBM5+DGQ2hk9wJMO
/IZRv8yXuPMtmbvEBoqB+vjR6POugdmAa6gkqB7FO6UuRVRbiOAsKwD/4VsXQtiYtgQj2+FmeoPm
PWRuSoZqWiut1BYKr2aZbkTBGxEcQgUZqUPAayWGiVlDqvHTH/jAA7KL3D4pSfaJRSCcQFZqnTBh
2LLL7U7CsSsWsHUEnbAoL0LbZYyIDEl8TBeCbcUEmF9jICIf6j8UAE+5oUYF828g5N+lJ2up6Y9B
iMwk6FJP7K++uhZ3xMzWg9eQB6H8ItLEqdUywRK6A/z8/7L73g83INZmUkFUIpKU44v00jkzJqyh
Wvl4dtKD9uZURURRnS2vwTnfwwAT25dNr80/jXvDMCcQqF0EPwGsMywHo+F8FN74k2TOZwfYR9JL
TNI2Zk/aG4R7z79Kcj7tKE+FEjiPNa/6ExtWttz80TuJp01nE5CiszIiAeNhxzrDDbGHrwcXleNr
tBrzDZMLtG0FvnxcOd2x23WqraIi5ng7YIr9+PMJhLbN8ETXTGniFrsEY6guE0mbgjX6uEMAPNxY
tfb89I+CSczS50WH8La4BpQE49JbA0VYu3WxasIsouNvh0/Stndr/6bg2HPgKSLZ6DQ28nix0lXh
fWATozBKP768mvIP4hzw3T0rzgcRJGJkCs2YbLLZ3U5OO3UzLLfEl+bkPPJ2xS4pK8yxR4J52gf0
Ma8RIwrwQkuYki8PXkVt0VilGA1pvyLrUgR+23y0sUqgZM4znv/fhQpcHGmSKPHTQCXjTkPUs+zG
bm85hdwaxPWGLMRyV/GzUWzUTQUZE78UdTtyBkhDnPGI5vVOPo8dHZADp0lkkiRDprHIDKq2cZue
xEi24Ksul8IFSpUqOq2u5T7oF+6LagJtSyo+gkvkepFiQomcTHCA8lXZKsbHoMg48aIgzyASAHk3
bydHTSg8XPON9wLPUqTG1bkT8fIfa3omdDDCkW6cNlkhUIz3G45q9Xs7/Sw50QGPOEjFIeZ+UlGo
wNAa1gd2NimyEcs3szUll9az1jlvW2tV3HBC8D2fw4BKaDdDnEdAEi28KzLSBWGh9fQFuijXfPKE
q7cyWk0BZWAwifC/HU/nnK8AERVcN+2vK0rowx8NeFx+7SCZJht3qw3RqFy06x/jwXup/Ss6d5Sn
t8hSfIWsSW05zghoF1xRK8h1A5PXQc6iqacicVTlF3XGkqKbx0o0pNNfkGe377FPm8zniNjBabT2
O+t2XLde/OyDgBHbFstU6iv67rYuPYIrdf9h9Q5eDu17uMOwlfsjHlUL4AF+Xhkxufm5naaLdhF6
KmY8sOct7RtxHjgeuYHS+T7h916hiM1YnpQgzQhalYC/LVk8lDROBp2J/p2L+UK4MGQJ543htrXE
ghJilpuB7EQDZtJSjdTKRRqdCUBYPxhx1CHFkUvJ3R/XRC/cBq9ivBbPhfm1gVUG2RyAnc9QJDFF
rYtME+1YpbNxM+w2cz/Z7z8vgvncw5iEiBEbojHHi1vCZg2GGOjjqtniwnaaaJkxdvVoEhlFxvCl
F1C2gT27k2sVC0zCKZypX50/6iBPaLPMleJTzr/OCxQaMc3AS60Y2fNQhKnunmaH6pjloSeoUV6z
nmiNTUnmOH6zf3JdnSeX8eoVMEg6KTrNhwhY/axrrCWkCP/N8ridG4VRs1H7crr5fCETYZkrW9+m
wo8PFNacShqjjyA1P2R8DCkFy3ntuUhCV0o30fgJl4DgkVRM+7H+hIJM/UT7Rw0RWmryTF0FBBVl
/4IKwOwum0joccLpDVMzG6I/BRYgWgzfIlfygaNwY4/F0yS8zvXyJZa2OKBFmFYSG0scJlIEL95Q
FRZA7nlAd++Rq0bBtylhl77c3llvokMHccy1Fkntf3TyCL3PhBNSHLuao4N9iOJzKjdjCU5pjPRE
8nU7GgbI9v9KlEmah2zbrzsIHZwO1mFxmyYj/NR/m/AR6ntSgILOZ7NyE1QZjniIW16LKg4+J61S
TupJDKV8Vmh7LBHPWqLwW1kmuomrbofJifcIn/MnQTiUL4AdsJ61d4JXWZJWmsmVGWl+7Si8P3lF
sseKE0XfX7a2Qxrdp4Mza7cX1TPfH+lTVoZOaQdlja4Ksqn0cS85c9PtNqrKSsPar7d+NQFpJCUf
pSHAir369d/6s7InpzUtNt3L5U57+XTEsAoWdcDicd4O3RRD3UJmO9s76vWnLWFpMZ/GD8opqC7d
ErKe73IIXb9k8HDrU9GlC8EiU+Y1V9U6etWP3XGRIL/3m2TsVxJKk9jIPO/Vn7765nh6dqoEFrr9
LOdo+yei5IU0yKcsuTF4FhlxufztLqxad6ovLsjH4bJsvd/gVk7F2Qn40MYaaphVK0fviTCa4iZj
r1VCO92OiPMbRAH3zgASRhzJ7O9PcCPYjvIaMCk1KMSZncyKKCm2q7SeUW+kQFcv0IPIhoDHcUIv
d8T6bVM9QGlBVhVkIBr2Lxxy+/O5OdZTGLEkbRuI1jdOO53lfaPTXLEJbMkPB06Yb4keCjik/U+i
tOnrF0NM29UR3pTsC2+PFgvad+Lnn1uiurHZ8ZKaUv+YQf3HOFwHgBKPS7KbubsCgtU5Cx91jRk0
Am3BRH2l3TsyfsIUzLsRh6K83VRSsvKPfTOCmqCnQvyv3uFxx09wBwyJti3xsOV/Tja49bxD/Obp
XUoVDs/APOZH2vBZSw/UjmohPQZw113j9RXUSbMonOKIF8XDyF5Eg2hr88NyojeUVyklHcJsUUtf
FiP6afzUOLMlf8g+JnmwkcBH+yBfn8UOkWFt9xBb7864abcGpAUxe6Pif9QyUJQHw0BB2nLDJhwL
AlItASncxpmUNxOzfym5iN4ZtagfalR6Rl5q1YinwCnvpwidrOloPlU1+FoVgXxM1sM2TEEVi25K
gVvf4XCnrLbwn8FobG1cF5LuAjcMwV539fDkokOOqZavIaRbIg8pRZQ3VoFXMH2nu1aGTjmjlagx
8cRLjDaleSq8InodVjAnkggSLT9b6DyeEVmhUZF9o0yeKTkLl8IWsRv/IrNKL9KcCcAS20n6x/Lp
/+iZTSAX1ZkXvaHsFE+0G2UP7fx7GrXXHmWtruvxFhzg0TefFEiCRkc3xnAMiS5AB4M+Fm74iFak
i02UKU/q0WiTmCLD1N5bc+HyH7o387j+zucnE/IgjH0fO4WJ2keDz18BN6hrmrES6gtZZ5mCPh+H
8P5S3x/st/BlCkfiJCedOy6kCdnS1RWFLe4uwl/iEWkJJzYjjqxrq54HLBz+s77b/v6KZwyOrrHF
sSHH6+U9wGdHPUHEYKBwHI7UmyzXYx3eajZwQFhxW+aI10Zs/zMJWC3uNDH1mmkMmws02hqr0DJi
RVfqBIc6bATXE59QJcfzWNALP5J8dOljueD1+P+wKw5SoyGPQ9b3PLmFDh1aLK9iirJspH5Gr2eG
j8vSlxp3cZpJR7lPPuIdoQi1VMlUYCCcHZ5iuowWh0hDwpz8cOUtPU8LuQv/7fGyg/1QPzQ5LiMC
mLrDIlblX042d5GybhhxtTHg4G05wwDktVCLIrNdTw/abpXAfKvh3x3rLsmPS0iVNjEKH43we/pt
xDXsR5SKmBqi5iUPX0x2WmfJsRPtSej7ocOY9OpL9Km4waoTibuALHhdygcLEFOMxuhbjjhKzS32
BsheVdCNnAv2bsClXP0HlHborpmLzETblk811xl0Cp6UZlSl/W4pxt+tmmjZqVbJjYlGfr7ZwuEY
8bGWN7m0rFAnCwaZ59hWAQ6DTPrafn5UFTgH1kjlvRSwiS59ntJM2uI/X6H6raVLbEQHoi9jtW5N
0W4GMFfeJ/qQG+/jJCFmooupqJiclaDWErhZnJGdKng12n+bGQvM4BCDFc42qzHRL+ePv4bCRVea
XiPUlBGxAa0O/u7IMSIxNBueIFy80Uz6l178Urlb0i7rd6zPAcEbbhH15Muq776WBhAoMO91zlf6
sYujrYxfaiZOZKMqqJFuzGJSFOFh8x4kvuLQNoKZdlDvJDAgsDEFAFo6+/skiaHt8qqaqxum1jaG
h9umCWNZQptqTdt+4ijIx5Ww4g9/G84H+dzKCKR8xHlleo1vVjk3MOLA8a/SzUthTk0kHgXaJKDa
VJ9eN9W0lnoaOKl0bKIq12Y+No+7uNzi3FQMId0c2VWv9UyeZ0lVEd4deWDrUIZeXr5o8qwIo1gA
pXxDR1LFuc65QssbBl2EGzSiBiSq1r8ZGREUqk6e/Uxik9DqQP/kwLhiFDGkk0gA0ekAHzIYhtYO
kN3Gl07QVS+cW//LYooFrpsE6Plt8aqmkl8+VnTAhMyhk2gYCj3t07rbkfpIReRzAAvTNeZ7XN9e
brL/19c3AJk9DTFbcXRqVlUvt1s/P/MqFT1oPDgEX/OC6sAuLvAzFpv8Vg8qjCcUqf6yA7x0S1a0
WWvKkWHcVvhwhiTTPDEVxMafYLjeiMmwoZfMjgVnVBvHwEw09AbI2HtcE2mVEQHbPMrUJsJA7K5t
c1xia+R52YivVjxU9kN9pLEku+71SzwXdtWBUTqUFIoIu4qXDOttHs3+OOvUyO6/RpDadPuhhrwQ
9qxEudeoCDsDyupz5B0aY4c8QRsjupY+yXmCYekHr0VQKVyJ22TfPokB2dQjtkQ0AHWNXd8jZsEZ
qoSRKmGjg+WwkI1+s4qwHAMHwV1TrYzD3kM3DK4+FdPO4kKb8LgkV01ozFrZx7svd2c8nn9+4M+6
OXfMMiCEpFg+af9HuksPoiBNU3oqapnrSdZpCaam53n/BYaDsokNPQAAI/D8rM/Bv0ZUhQJe53Ev
5XdDdmk+NOPXxQ0LJ+fkVwpHLjlPyLPgxF+1N0beUJwESGfla4lM4Bl/cnflrLscVYJXg6Wvj1Xk
yxmPR25s8y4Lq7H3oSyphz6deaFiLRsKC/XNopqYuzHWcvu/FUmohAntk6BTd8kPmSlpBTSAaKoQ
kEeFAdRTsAXViqJotRAh2JbtehY0ILrg6DaDQKQ93BvxTUtP7GQJGN5R7gFn7uYa+w4rxWTbc6KU
xpL/HZjYt0L/2fd++SpfwU3Ea6zrGSafbCkTjTLE+cKP/+6Ok9Bj9ufdf/kAhklIN6G2RPhKWf7D
P4uSfUF5u06CZAIUIa3VUTzlTBXjXzQIC0OmIUsyhCFkf3QVw5MRaKHujjUm/ajt3PEl8/F1zyvS
MRqZf45HuZq5v0XJbpag4jUjIzJaKKd3AW2Hmh1tqcN6iKYSIYIQQWx5KGZeev3N0PHNedBVMQzk
olx74CEQiAdWD0UmH8N9MlMi9zpkMdjF7mcBjb3KMv7cGjckAAOHbsb0WHKkVMQSBjnK7aZ6dY2x
nKfy909EGOoI6rw9pHUJ2Dyib+qS2EtOxPG1ZRamgFf8qM8B9NNUz+csjPiOlxJvPOFqR2elP9vs
CKbm/AASnVJdgbpmcWJVBj2zYO829qvMoNYheofaGVNXNsuPL/Qug7P9O7Z9Ve6LwrpREPYlZuOJ
2b8V8WXZkw2gn6oItXSws462p4XccLE/6NJ8LAqAtJFax4KGNWmcO+gsySEWC55A3HHLVJS7S92H
Lhk8tOqtCqiPS75FRau3fE3o6v5MOg4TF9PPmLi0ondv+ZwIteh/ALS+D/nyYMnUrD3iQaDs5XOs
q8JCGYsTNhXHbD/FGeg3jO+FsuaN76z1K9ZMD6861vy48JtmAFNuu0j1c/2e1UIboMU8C/NMBj+g
BT9qusbDTH36fbkK6oe8Vi8HG51tQFRBMdFV7LTZjOPUA46N6RySIUBp8voaeVvOMT+LRhvzwWm1
d0+yTquYVZLYSip0lviVVbdY6QBXium1L6eQ8ARVZgaSYpQOokaDZPtiOmsSQpmCHVpf1sKr+L3V
gV6bvSkC7kZNt9HYRlDmTnW32ViNUPXKhqjmdoFTy6z32S4YFfQTWXslYlSwGwnYhf9YhCXsaKaZ
WPu4z/KJM9KIzFP4u1XlTjJ6aNRsa+FVYjwoffgr+mfgpB3DmQiaqGyPf1QBmMB05vKlwmSUPSps
cexL8VDXC8iaY8ywCvvemWqmgZHmNlQsy91UjM21LuKFcrPIxhRefRwdn/lv/DKjM8sZ5kfxaIIh
98PzmGyCiu2Kq7rm94jA7o5FAsxo1hEbC3BD4MVubnDjGH6v4tWMvSpBGQGGu4AN+f8hn4Qs1DLp
JzWzvNAbl6i9o0P0LXR7MWCVV6uzomft9/zuoD46BQOj/oOmwokQnjtHlvQTxz4qzD3hatyvUOD2
/5fR/ov7HZgTyILqJbNmzwNUBCTJLGiNc1tD53oY96QfuPQGdUiGCqEPUEla6qfUe5jh2iv0jbse
5PAhQagjr/XgbIRzf77w46qryjIGKQVw2sKZFgtxkSfrdAum7OjC07vNUgHpW2xZCVpLwIHhOBUj
P7ExSAdGbWp/woofTrop286LjkoT9m2tw5CMBitUfQlg99JCsEiCazudDFIZIUvrp2q/CnpF0+ln
FdgwKIzZ7SlRNmFFDZcY5Epi9v/35OzUxiCStGmU4uvJ1/VBlIkd5uQZsBgMF0Ja5cIgU2BQ+eU+
0+GINwiFE74vyO17xRR26mx+OliR565TKj24UF03zqezM9hZApERqjWbsW6jADCBPCVEIS5EeclC
0qUyIX2JicD/4aH6RsoImKBdH8LoPdT5Bt1AS0Picg/L317J0LU2fzi8iDHkxtntpqFpltx6/O1H
L7N9clbDed4kt0wV2LAAhGRgwYnSsUo9kvGXqsLjTLWDC5T/ofe6TqcAC1tqS5++h6/O0xp8EFyM
kf+Oc4Y5VHJj+ZYpoX9zXO5qgYKe0i2Y7vkYewNw+6hiwVuS2C1m4pJSG2L74UQG303HBPdQ1eLz
+XJtA6m4Qkn5Nqw1ljupDYJXwD2Is6M2mFmZ4zwacGkYp70Q9bKir5b5N0P9y+ywGTphL5EMaJYT
M2WIt+710jQnN8fC2KK+iUKt2ps9HdjVx/V6p4hhrJnf35fORKqZGbmuKFe96ROT1mHLCx24HR6j
BHieNWeE6GBErj8DanGoKCIZASmJ7k5LlHwxnWaZtZBXJPR2iPzVlXfBY9jxreXBGsKkazPxBN3d
vTwBbz0VHHw3h8MRdzohrWKLk1QPUjnh2CGkqDLTad5hUB+a8rdEOSQVN/Lf9DR/HyrCGukXYwJL
UCGxwRsNh5iwAi8g76YygwLDlecEFOudRxjiqZrd31vbbr39iP9l+PnOSBwjFKNfsY1zyNZhe8gt
lBWXlnhYXqa5I4aWDHq8OqctymvJ1A9cPef7FaPaszs5G4AZzuP+mFjyxemeWarZzaVTcQ9ATyhR
7NDzzGRcQq5egH3WTMIEyXGORAScD+29f+g7M8gwjhM3W50lj9/JFy+EBoSZ/9W6sGllouBPFbHF
zMT600qFgUD3hp6kQQ89nYPcc9CUR0Ar3Dc+bHT/0HVG8noYFJDJsV68eqIW1dkt5epjLw5FnSnN
TroRH+I3BTG8SkhQKexi9Ci/iRK6R2yOBA9NJv7KmG4PXkRS+OXRt+r84S5aD+rmRwOLAr/Mjamj
BUtWYE+uHSb7DyG/aYw/rSQMLpjl607nhBwvK1sKCNSS/z8nIoktLktCkVSSS+0fxDHkv4kZlSea
KUtWJlSj+I7a9JSwfK6QuSDQ1EOL81SvaN/4SBn28x40pXpFGFSvxeUaBF+V2P8G7cT3SUPHdv28
swL4QGyZyeD8gZM70G/hRdlNDP0OrHn3fZuGDcOz0RfPels9TByzrZbOEuiXUF7icDATBLRAVyK3
ypse7EKoKSZ3dQBzXi+b1YNLz+Ooorj73LT63ZJLloMjoXJP1yoO2o/x/o4dBCmwTW3GcIQkIbIv
Awz3YRcCcFRkYfWM3KvqBiCCQvCEwr8DuHZkRsjmQkEx1Es7Ee/OtrsDboxdYPD/Km38PAaC113o
BV8t85nagxYiuhlXgbjLhvkK1Q0mqpvIrVF9da2glb3yy+F2H1AvGxmaZtzgbOEQFr5TFswVYCWk
g66M5g/fB8zI/mzzOYXbKjEdcyCvEtP9JVN6hKIozG1X4a927fgPfz8LEQBLSIMAoZOWQEsGcKFn
bkc8VDjZvivbs1BKciJiP+AjpFYfbpanzrmrCyPOZZj/Is0F6fuyvK4oeB5GYlNOe+JruMhFKbYn
eKSE6D01j0n/1lCx6Bw4Mlb864r/8qGFy8DFOgFwoFQbtODHDujtvHI0u1jk12xbZn5uTR6yOPoT
PYNgYXLKPYi/aKlOk04VuVVY+53uR3UOE+DWFPv06g9zC0HngYz+O4g7mG6M5IG7HanxLVchkDu3
/M/GoHnSEAxEl8Z2wfygUbb8KQcEVkBfXctRI9WpDy/fHyO0Q4iEpkQM0KkPTazK3dbAMUFNmo7m
oI0J+9+CpDHUFXiIimyDKYfFGqkMZ+BpZTyTwZmmBp4INP2OHA9srsuyQgVFPxGc7BwXN/PJqW1a
qQp6jtyxwiq3fOy4DO9iqpYjM686sdMTeeVkki1P89+4KUPGqH3kBv/nJIhNpy3eFhjCYLEFY+xg
ZwsCE8V3tTQHyUaPGe2+1IiWHOAsQ5xxmfRd3Mx+Lr1Zp99YephQ596NGvzTNQi4Xjj4DUSItR1n
dz6AOsovthepbL3au1tAzcb7hLQROCO7YQXU7dGkvmuYYqM7I+9Ad262pOdTzNRNXSr2rhYZscO2
KJ//IiZAVcWcq8m2e8EuspTwYVYP3NtlXv16u6q6cAlVIaAIuGynrfNZXMDtOqC39kMGNMqhw7O9
B+Zz3O1VtJHKTWP4yBm68h5OL6tbya/dBYeAlzhmly3Jaofw2BU389pIShGtaKoNXyLv7kP9eGqt
1iPpDqBI4Qn6iA8MlhbP9Xi/pQe0EdLEfOS+OjSLKR4hJTAuOzHqNbciGWLFQkdkHVfkcD54wEh0
+TicZ2DWQk7e0qD2RJNEaqC+RUxGpXu5dQ6zw4JupSRGMIm9cqTB5W75fFvppY7E7U4D1FGt9TtM
Dw5D2wT6Q6XgBSwy909wscwRN8tS7pXDtpS58DuqLPeKUWWXLORPblrdlk/0LaE93kpIxFV1aMn2
BObTib2qdS6+nXWixmVeI22izFiRg3SlMz2/YnxM7G/QC60uu3/+a9fpTPB2UQ+oW/D5G8tGzl7C
ceguPhT2+cUGQkcjGEx9wGOwJB2dq/S0aCUHDwypazH4MkZU7Jk5XNLiXgxZ1r0bnyUmQDafz5Gm
6hDuiqQ4q71wZSQ+VrCFBEL7cOhwBBAkKANmIfscI72Ek32RDpflXKP2YecuF/OPwfgfyHX5mIZg
cpJEBmlijJCw4O7SNWtjFHoEJ6WPRAnvg+lrJbqKmf5ozL64yY2rU5Dwiq8ZQ1znhMit0XYbqUli
qNF+2j8V88QNpQ9hOQJvf9la6eUyh5SHjbEaQaGnfEJI3Ygv3hcbpWndrZ85itEjHILf4pitEoBB
3blGalrMvng2IGvLB2y0tAiv7Jyc+wjnzbmY/IpURAA20yQlsS2YAu6Dc45QHJxGa/atvQZyipQZ
dMT9E9f4dhOgC2YdA3490J4y5uOAXdhKQaIcrXd9o9yh90fAddSdcT9pzujU0NUjInIM1ovo8ZfN
F5pAb+papCePQLsw4UpW5xeoaQynv4O80/XFvmNq58BmCgVnuWz5IEQf2Hi5TM6TDF1sEBXUAstE
f0M9H5GVXPObmu4pyYL9hJcfbv/Q3/8QG5QP1c9kvXAz2CbH8/I6jF431GTjWH20QdI0GZi22IJB
BwEmlkm5hgkbg2QKxOemJ0L9KgumrVFb3yXd0jFbM54C/EmteIJhSGsXd3TObfLJ2r9mntq8DJK7
kllsNZ3jKHxDJ5wVOKhqdgJ/6xBkkXUC4+dl+ee0YDTMvHd4l+3gpKfyyGgRn9aVZ6lm5Myd4DrP
xsR2KYWFJpzuz0pg+cVw66h+TI3M76aq8jb2qqvngGU9GvD4jUmYGOOWMb+UZwwLvELrWyla1Usn
fjrJCdDrNKbs8PeSzKvaucP4LTQEhQYgwMcL7+R5Tzre79yBEPIHzuDgBeDygtly2Wsp9c9x0lXC
y5n0Zosjw1SIDacIxr0bwqkfPfDjCDQX92LW65KAyi8V/BoCMa0igS06x8wYKAIm1TKwwxGktox4
mrFcqGkZaFcZQRK1umBAYm7vcAcTrb9JJjOGxkv5Rv+xVVA03LcHD5eBOjFoB5umWSxh2kjCop9p
IFQLjov/PqBLdY11NmB12iCqVMu2daJyxEysGRtziByAjdupkC+Y8THr+pXZkt/bxsNreFLUGbU8
SHcsynol4KJWod6W3uOQXJNmDTxnaIWmM6P7y9YgxkI6yEQCqMh3yPaar7Lk3YHmihxA9a7/qWMq
RA2F9ciEGFmsy0IemaYG7QeZnKlkggaD7R28FXjOkKJe5c3INjH+FUBWWR28kFZd1euXtpHy12a4
rwL3BCQQmNy9yJnqar5P6qs3SmrURnrOtWrzG5tM8zLY5FWEU6XOBt9LThTIlSrwTdtYV8glrmwx
oDvwu4Tb6V0oyNCO/6IzVN9S2oNJXQeztsdid6AW0GJzzOhMxJLIUcZsvBOJGrTkXjik51Lfl/Mt
VH6aqjSUuLNbNqv6uMF4ByMiD7oEMAIIwQc0i4tocZe4ZZay0ZgaV7hiURBqKk/WXv825EEh5dcC
PcbqVPSDRmoz8jHtIFSyAUuqVshZFQUIS1qVyeV2d5hhg8bypJTQj2mx1e9pBxJKe+VI+3G3j9i+
q7H4jH+6JeMcZOeofHU/kYoWEnt6ai96eSRqANmARUT1HCLBHBjhDba7DRc+q1n08R1/9JBWebko
oigLy2pIGf2p3jlsA0Pz4Xc9DDjyLe00Z+Duk9unAuNXPgeGraNm8nk8ThBJQT4Ha2wExbaHrHL2
Kbxjc5O99o0LsHA2UX/Oe26HDS7gGLfF56VJQl4KCf7zlkgKnkhksIKsviTbtNZwm8agTPCsqcax
rAXAZFAisb/KonNxMMBBE1Zek9CV6Tj+SuLPfmAYZfrJYFUWEne4//zZBtKqTzTb9kYfADpOfH5f
Iv1UwzP1vnRCjAdM+EFuFYIp712iVrfjCs+GvpW9onBRUhq3BFxDINQ73O4YgqMCmriSHPRrVCY2
N0llBBzcAwFDtwAFD7q9hPGKoCzRPYvQbEHLP5pZE+Ywq+aGp3wEMw9F1ATd0WNgJ3QXoAIZ0TxR
VgQM4wPvi3MP4gt37+Hh2FUnqTf8MZAeY2USyD+xvp8X0XPOguGxWN9UkbIg9pWAnOlW6oQfQRuy
WCdO7gOGuPfxUQ9ga3X3LEEALHNyipHNEDFhzkb9MJWZyp7jy7rEnhifYs7gGAL3dlSh+K0xhGk3
enM90DDmxg9qzcH0BOvOXv4bFRixlg0W0pzV65aQS+K1lbfKAK2X+rqf1MOyYIugvX5GSWINONQa
ytLQARGZfbrYuYhYhSUcIK5vULdjCJ/hlz7f52Q4yNHDDzREGVfcQxhWAr5sPyINlH+w9w/FhtX6
3N48QM99zyoulqb+aaCC8urL41VQ8cbuzdkhuN0ipIyGz69Isk0DojMhif2pSAiH9i3bokll8UYn
UYfA7fliQvtVQLs45+RMExKvrgIbIFlgHg9T4A805SZtGQfFcPFZ+njA2TjRWdKJkVaXjSHH0nl+
M99+0sHvFmhGUCoI7HRF+tUUOFF4djSpwPWe1sUB18SDvWg6kfXa5jxS/EY+HNZ/35KDIDLNDazl
SYW6i62CpfZ71cU+xua4CWTmf29BGrPIesfS9UL+NNVtAMvglNVqb6q3UlpTHkHNas4jLx8PZ8+5
9Xs9qus//niJJqbu6IENFGQSEAkuf4FqY6OMB44xv8DUT4doQ67PM5rG96a2/3t/MFYjWlBRKsk2
XBpYW8gj37iobXNTjcUBjHAhpldzBvM95MbUOw1RdjHc3cvCJ0gTeZVhqhgEE0Kf0uGlfk08CKKE
6h+1eytVLXDeao/1kvMlzPk9gHgoVpUq2/AQenZZ/jDgGvwc1Ymo5V/LxXAvQ6AcjKIcTsA0f1v5
1dFQPUMIkqVHZuKc2gXFUY99RgcEHvkE2sJs3m8gdDNlA62V0nOJGEk0T5IikvwNyfpcaH2rz/ve
2ygDsFRD7B7qHqMDNiXkH+VZPWSXHom3KKOXE3DUUdcf+1+CP1APfEIp7JComy1Rr7qpfGceZ6iT
uO0gMA2QQErH2yjRKqc4784nkzYMdoJ17A+xtkOCGlaFpLBL2B0cdtPEXvcK0RK2zdhICd5VinfH
TsYh8zWQ1vN6bNrImgNmQ2VVNKBzIq0PYnRYbOUq1q8SEnZVtqw3n2cj0PsxwfYkFceR7NwcAbMG
yUHZ4ZMkHEVDKtYYEU5weRwUVeMX5eogGa2CWTD7Ml9/eEEBg43LxYaIH1Y7yhZj94PMKN7icpLm
3Up4MGeYkz7xZn2bKl2+ui5N3ICCwMOlEtVVeKYI3N5CJQBVDMWy/GipMgHyL8J/bPlq5nn6jrxt
ApBjAJPJorHJI64Vv9gYKsqtXsHkIZuS5yDBemj6pxoGrKGQ8Wq0TijVuWT6EpJOfpcu1XkWRE37
z3V8VI8KPB9eQCLpYOn8FMeKq/BcSJtKk5kdAy6Oj0l0AZlVClBIHWR2odF1AyC8VRnV4D8LFcl5
tR33RELnjR3DP738JAMA/+KeLzDhvcXr0l6HSWaqgZXEGDkfAgkzy+JM+MvECWYJX55Zn35YM+gt
XAGeZhthq9IUtzcGPEcB2D4Kpsr1I0IHfMFlg2BEnUNdwy4T9eWCo4sIaZZvpuX/vvSHZAkWNwMz
q9xq511Inv4NflRbviUXb7ssW+kkZFperXQKfn2veD7qArZD/wxllg37ELgqBU1XYID7vYQmdaio
ViI6XSNsrJdrBnObRYuM9UbJ8ZxMfQeI9GEanKFaxxTJwc+93zok0Wo/4z5b5tEbIdrQmPAFpG0G
aAl12RP+YIpx0wVcsYWQIXvIhch7X/opIzyDIYcoKzmPbTISiiYrtYhldKcCcb1RLPeo1LF/kM7h
PSsEycaVT6uTjLK6iSxsUaeWdvXQEycTdLwWtBlj6h8mkeSbY0cmRF2tzAE3Lr+mCkA5SlseJ9ob
6ioT1ixdu0p9FRb1UVArsQ06oCaWPtGDLetFG2MSucRP1B71tH++cpDM0tBLuoiKfwyxFqSlG/in
76i+sRiBMlsa+zUh9WvkbVB5seKmbnh796JJypHTGA57pVB3dTuHcJJVj2dZ0OpR8PfMOGxlAKnE
vKI03nenK1RQ33+35wQN1uYvI63tPC4IV52yYMSx/PG7s0l75C1SL4ALxnke/lohxiG7ItaVt/sn
8pfkhsaPP+KM+I5bi2mQ54nYJMHhFY/6OML5RC+CWC9oj4gTpZdChS4k8p2kC8j31EBrR0flXACk
ovX9PmLKhhB7j12poxAUFvhjSl5aCPVhoazXaM9aMHtsibh61I5gFCXwhDiKWsGWU0vh3Dmh1O7t
TI+eCaAt/SDTWDRqLoZq4wLqJkFBO4+O5h5A5fe8tJqdY77UR1vr7JyW34si09N3vGoXvnuSMVeD
fS2ukmwdO13L/v7nl5XoHlLy4MBvTIk+Wgdu+JZo6TTAqDS6t4PHNAglJ61SBvj2ikGZyheLyJZk
1ahRAnZqQHvlj+WJSHi467MljbaofZhKJdn4fpGdWhDx2aK+Fzc9Q0HcgZcCQDS4T9hQspQfzs9E
xOK87u5DdtgUnuVO8R94SGoWPJLoknB+nET4MS4MRaHl2uwo5CtNLUYPvONZFdQ4Y2mivqgAfT6k
DvwfZ9tA1DOw/OWhRhVXu4TcxvKk5vB3pNF28xtHjnzQqHHvwC4vxonmolo7kba+9q5iB7v36YNj
wslz+O8DFgXSHdgkmxCBd/xbBQd+iKD59CDRim8ir9B++IG79Iiymwl7JQGwZ3AJ/K9lhXlC5Rps
p2djF24I5Vr7ss+EfCCK64WSUlLXIlJh/k82cFaWQKnoa9GnytFSQzBq0vmhehgfqAaAn6ziqs5T
2jz/kcRAKBToS1/SLIofxkTKxGEPFJ7T4bIX61YReizpCf62FGL3nT4QsktSnl1XA6/p1jdPEWNE
W5cnYgK/VV9htXAgSN0H1YiAK0emzJLdTgeX+AluE1uSfTzShu5wAcYvwBr5JeUpZlfA9R+SKjMl
8VUOkkE5fZ/YeyzfQTFSNA8tRIgxcNd/reCPVcC+9spbJDB1G7EvWAHVp1sYC59LFjwggbHJoIBI
zVVOXwl0/3NBLB9V5GOIItAypDfq9ECJ9E1XxXZ4ZZeaMYt0seK21EWsk3XRH1u7YSwEjgcYghIy
Kgcw8j8ATYn/VXYwDIjP4IbAw5aRCcnE2eUtpxKjr58zEE3WWL8Y4wGbluprrlHBJhvAiEVrv1Ga
sLZch3qJtDezNxhEZ7uY9zup5pSUzk3k8EF/Yg+20sFpZdzrNHtZy2QEtQTTsHQbP9Mr760vP50C
Hm2e4tayr0s6HpDwJeJY5dTaco6ODWHQ2wXHNjT2RuMzyE3UjQPXu/Js0OqxAiPQ60oZGGLiVOAy
pI9IxQnGEdvA1CTx/W6COGncIb2IrHsnTjlNtilxSa8OL1kM3vYuAuzzxVYJvAlvlib5H9YVv3+K
cptix5pUEX35dYNwADjoGEHskv0NUrhGmOX6NK4ODSwJZ3J8dSyQO6SZqMRZbIoGwHJoco7hr9uO
CfYQxiw6FOyM3ylDnj7E4pEnL7zaAw25yG2isiiMerDWAYByI53xqBFTXb3VqE9wN64idsHQCxs/
sxF5eU6bOTxsIitLbiZwgpBkyNQzzku5BvsgBLC+yeqaqRhOBgvGK0N2aYDmGg85PjO2PxOqTkn6
+khCihNGVQOlY85VCxC60SZng8idMuqf33+EaTMInk9ExfwT/hEzZ73S7FYY0lWM4uN/axiCP9M4
8hORGn2TqYk3W6PlwdI0EIaE+sLSkj8GzQnfVuWpbV7+g0QyOoG7zkUJ48yJwGtCav03zHGZBmLH
gFJxLV5k5kWALTbOKnWyPCVRA6zf8qzlft+YE6HrP7F7slF0jFZQZFpXPUWYE/vPLZNCOujIIMid
g4dFNGcDjaxUezUo0HMhh/y2fmFyoG1T+GRl7/rwiXceIUxEDXN/oZqNOIh9QnA+9GjGcEyX0u4c
RyOwAnckfy6Dl8YZYQiSwYxilQVJnofZ9RC1o2gKRem6gPpSDKeuJ6VaG98xbuF/3CmpV7ZWyXEx
rrqGavvqGuD351BVvaw9GGRaSpOwfKa/CDAW5c/za1y2IvDYOM47CGR3RVYkmxampgR/irpLon4B
eYT5kRXzLUxHOPScbY7Haamj9mtIKaJz3TjYIfqu0owYJ/HkRvW2EIlZjo8olTprSM5Rw+vPh2Zl
aXKD+JP0A7WO+mNNuK7p6myCwtLi14ha3W8e1B+LmrzdyVBHaIlC0DuWltYOrY6qQQGPDA4nxR1n
Kw/MmetvMP6HG/V+nLw4dLdhKakCDtB2xT5xnUEAxN2GgQbaEC/XbOIhiiW/WXSZtsPmblfa6zFf
BC1nHntAJTPM6/YDGugSGJaWxmKgSqVxQ+zJDrMjDSrR5I62jNQa06yhmtq3bapGU7oVqTYSr303
KfoyVlt5O1Jvi+DMueXJW/n8UD7FpzDxXbjTlHytbS4g2yuU3WBZu6c+YM8kfrgUWoxPJcx/tUNl
t4FEZUVK5HYwQaxk3CABpV0tml/luueyjyxKyRbv/a4GhvvxO8K1+XAeGc9w/AplUFQt5+B5vGFY
EYb5QQSCFJBtVNnq767qiPqt6wU3hNEVKbdhfAuIkDOYDPH32JCmNT8/FHISYVwnEVr5kSYjYrub
ep6JtdL7R86iW+Du1Z78d1MqOrjjcZcG91RyNrGA3czWKvAVzC7kQ6l7KLmfADUfE1/maGMH9Z1M
pXCUbnsCByW2XwBYF3Ho7v9SJOvm6XnaRzfYew6VKTVSK/RxsWYLD4sja/D+GTZ2rlwMSoafIgfh
PUVabhXB+hcwfnBCyGdRWE0nFCThaITJ+7RSqUUIkhQS73U980BKO6uo8DJni0NV8N9Xk5ZjJGc3
r/AznJy+djqp8kOg1rapi1b102oRkskLf0MSfGIlO5KhVP5ZepAU/obhrdrH+mRKAV9HsKnvfKWr
b1ubCKLlFpV6KKlPjl2sPeP/LHCVWhu53G9ka8+Lpgrb22/90QSFyTEvzpMwSUkYDI1c6lKnlz7e
HfwrqPG5/DW4wesehe+9q+k2+DE5G1AIpaslPNd8EfZ4gDdWwdzloyc47dFeyiFCBfj1Kg4iY/ju
sDtyt9pjPVhTRhMFLYEcwvkN4knKxzq3rfCJAuDQR7GAzu1qbHgUByoUt+XapezESDuAXmJ9JIGr
4ZGbFNTfeQ/K8TcGuekzxe5GWIKpN90fdBfigIqMfqa+JRSN+tNJ0jEWXgVAyuU6iK5cbtLCVpfm
2/d1qufb6uIh4ujsM5oxRnwtP68GhxV/cZUuCvVHaXE3I/DJpfG6ltegZ/8FvN7DCWEvHeb4uskC
oa5iqucDEQzJJh56PTo1Mo/ThpWB5rm7vGeSmexzmVLsmLzrNo982UpXyLalKn8SsGux38NVF3im
P39dQ8e3v/VOmb/6N2Ay0+C6j/IPFFwGWt34Jq0UJ5R1Hxdqu+DcGo28dn8pNpNLsIvCKTK2BdJp
1zt7j0oCl1X+vOwYMue8r+kKE/eVyvQ/80UZOs+SwV7FGOCFgzvjG1l1NMV08fY4bbNDP5/g682v
JdwHU/p7zHVIJImorYvAUIusm1b0O2ebFCAmOKRfyMQwksJ4iriO2UAN8zMw9pkqJgD3pNzozE5I
5nGmcQdHcSmbgojaKt9LY/huY1wMx7eBwccQfwq1GOQC89POchVSr4ujs9K/LCcnmVqXzplwQosd
gRQUtkvlLc4c3Ays3sq7gG7MCluco1YZDIJcvF9akHQu8pxw3STgp+ql2dMrkKZGGU2itzywZcmu
11g9In3KR8uxpxyIzbpCQt6WupFAmMtdQXEC0NEZOgZN0YRtdNiZS45IFBaFeLH6DDy8tjLPm4JP
tSGi/MOL8X+sIwdxIgA3EN5jHExgspMLbTBTRbPzbeJgeF/q76J4De82F55TV62nybcZwl8hqJO1
OF+HUrg3hVoiI4N1m+X4PHRkLNcT4koSyv3hWzeTkUyz/o7nyz+6ObwdwvfMIf9+E/Fvks4XDS8u
4qtMM3+4eASwNBT8JvPgzpkKDQKErT9n/AmK84jp/JxfcSp/ZjThRxFlaB90vV1wn32SQxuwTtRQ
mPIz5c4edKKnUvcg2sq6klP9t2JX8fdWvwxvzV1yY7P9CnmhrFn4nPgdRzMpwAKdORotBykyXora
8Ozti5GSIL3TxlH/SyzjK9N1BkBOvWGAknOOvpJOAhpI5UcV8sj8SZjca+HNJOiX2GwjEnIXeDEg
hsHZme22FiUUhL4HLT6Ac9PIw3hbxETgkD94sot4XhJFkAFHDqCt0p4OnUdMmWljJlsuvqTpD5Sp
l1x2LrFWbW7BNrp2CTaZN+KrmWcOkpKEoDUvPSsyQWffXXdftEeJK2e4m+ty80ifwYrEPDtk90UY
RBGfXA6iQDzwu0qHYSXf99ZKYGB35bjM/z0enFOg9S1yOWPbba1B0+JpcVXc2WvYhMvIJELTQrVC
N4H8T9IAhoeEeHSehAKwMBN1OoZeon+hoJbHhgCFJwfY/R7Zo9SDwgzWlkEVdWpZrpI57Fm6SUVX
ZogBklhTJDPVJg6jyHpjuhVu3EILJLL29UWO8oR6FHTmNHBrDFR2DJkH5iVIDS/F217H4Vy6w6hD
rkldaIoFsAMwI3nUUwm1y05ELEf9pAyy/f8rLt3xwlW2YbPI/26uFrctOhy2AzJvxS792Dv3DlCJ
3AdNOGPFhSpK2ERztI5M3VPv2NJ7CwK79psF+WGdvHbfEZUd4LRdpm4Jv1X0+8+8nqhXGj4Wd7xl
b47wYEWsB161ZaKYfUlYuGDzqQY1S+9ONJjpxhwR39MML1f3c0arlQ5IApeexIUp/u1PITolyRRm
x/+5tWprpuxcr+Dk5xzJrz+mWq2ZUIht4cmIg1al+8vwyqAwtHvx8jGF7fgmgvZwNTQ/vYJbnuK+
o+8cjE8ds8ywalatE1uFt7E35jMa8JGy/fJiQoBP7QW374TVts9o/kmm3+EFPOWJhZ0xVgduVxka
rBBrLjD/g0T6A3yT2LtO2Zq1ZWFzVrwvrmT7sRYJGHnQxFKS3NcKvzUUH5V0/tJ128xm88SDatz6
cXM5pHbKp94JUvo1kuu3Z4hn+fiumKX8I+NCBcGxDT+LvpW0Osa8O2eEnWQkbi9y5GYwSITKwyOV
6NLDj7hI2IkuXvobGEi46YyWzp2J1W2zVrzuHZl2WoKv08b0PTmN+7czY6IK4HPkujzzwvEuVUXG
7m8CMfAAvNHiNaaFx/Ui4xBPByAwasrKfQFEji3MrEHYzVFWuqJYqhvq/jAMrgSROEI5VFxHeUUj
HIsmEuRD61ARHgGpIm6E24VN7WHZD5noTKS/bdyOq30+wiL+dqGlatmX2p2awMNVMXMDYSt1mJ+6
WZPk9kzd1YxNMdR+Hk007tGT2L7angjgTR/XuNTK/AAjaMeV0ofLV2mHm5PLUlU3glH4K6Nvx20M
GztpXapFVNLnE71H0GHy8KiWsm6DtFBMevpZ/aVw+0B3HExSjq12kjAnm4S5SAwWeejZVPHktdhi
isGv7rGLX2botuLHvyZZjAg1LEWbsOdEzEWqunJT1L1cYnrI4HgCXXddGwi3GkUAJm/G5zsVaPA0
TQ1e9+jkb0LU5bH8RqBS5K9GM1/6WYB7lGWRS1kwxZ4QSn2n7hCMazsNpx2Yu+D8ISVtlDDDpmE/
J+2EHbQ5D0TeHA7dt8qi2htfVwdQCW6z+ggLYWvb7YHkovlIIrNQWofK/zbVSsDdYXx6L+FXxeOH
aHIm76QcDPmcBluZ9JaywweyfFQbbb25Ncqpo7N/bwjEl8mRmV0DTlBJXokO9PI7N3xFbOXtAT4Z
ajUMZxY1hQ0djXJuF5y3XpubosWtxVcOBWUR66Xyuo3mfI/odxv+0QlRfxbCsQ2QX7i5FTh1yxJV
JvF1Q8Tp/x88/6SVFZrjX4qYZSMXzwqthf2gTHe+S2e8815zIUEBiDz2QERR6zF97ZcJs0oRA2mD
Ka/Wwjh6FlA4Yq2GrMdfukdTD9mVIOszTrXXyT7517D4MQkku+vKcSgXR8UMmY8ihgVz6BMj3H7w
dcHaE3L3GR8+IoReb1bu5pjwJepgKoCEJyr2jUXMvwUTLkDE8W3BeDBHymjJHM3BpJvPdU6KHW/H
OBkgFDwFyhGcLED+6uxum9ZFxH8uZmabSDf4MyFka3AeYYltIC3NqleZmZkqFXCfsNQaj5ADoLTn
MXVBfSgSEfBVzWeyNvDKNUiW9gvSsh7wu8qgLMbITw72w/P/8rk6Q/WfKDxYnXarLrxBjZw8rfe7
1tNIs5zWKYGot+b1ZVXcwTmZSG/P5hFAjr5ohztkKX7aRmmyKDbe/hexp434FSIuGSlrskTUkU1Z
osfYV/Uanohc6YGEldUUV0E76DUiAYdIsQHANoHA7oFjWirYmoDIzGPfGBHHtE3tpTqK2nfRpUlx
HL3d7KS6WyJ1laiT8+P8LEm8yx+jtRwSJokBiiAdq7cCDu1hbgw1fvZVTbyMt1dPjVQBqvEj96fs
pQi7QKPOE900fphQqyu/f6cvUJiusTgil1KnKwHlKARrAjaUFWsuMgYF3QiiHY/61v7e3ImX0XJ0
pZDGCS72ZZE/IIzQk2/EIP2vyHJVmBcADQKloXsdRLBzvQLLt3xq+xIySeM0mbpmzwh9EdE1yYsf
8Ab58/UwpYR5mJucb88PlB8roOoN9gxaWXQkd7iPZjxzI4Gdp8Qee1O+Mr0DUhbBX8Yuw91bWRDP
2P2tOBW/3tIQ3cyaQj8X5DowdV4tWQ1POB/OPqwCPQ3gO/HfSGbHagxqT1/OwNcjlOmT2cePofM1
AppjFCkSs+0oW70UKn+vqjqdITzkyNmD6PtfTR5ZVCmE+d8mgiBYb4/wrLlsqNItzcSwzQXSh7Hn
Frl1ZChZ91LM2lAQ3TaAYpcZ0zhXhtoQpLKiRw13nbXa1bXwjMgOFAmzzoDnEh7d/N2Dtyqpuh/C
3PXKdTMOn0bNJjN/K3/z0G2Pa+o+eOpo8T3yOPHrnGCFkf7O10GWkWxLdvrnHXGf2a9dpuIkQ5J8
RJOJpboeHa5917eiwxefLqzGcbkafVVXZDQZlbvXCPON2BxQ2BPaNH12sZ0SIY0Q7Fx1xtKJP96Q
mXDFKPwllSMY0OGdZS3EgrsOA9pKxDjgvKyuMu00F8dFlUAAwSQF5CIREHmyRp85aK4v+xfS3pI3
rwUYF90QJ9vJc9fY3Xfps9fI4b0nbe6tyYQGrT8l8UgBkok/nUy+4Kvxg+lTc44ShWsoSxrj61tC
+POS3r/Ciwwplbx57ZkaS6t83Nn6ehTflnJcIxP/BVvsls7nhM+ayPXy2AHbzD38D3NjBDDu874F
8CqK7kWlswzjnbeXGAwgS/YuOy9rsLy6jAcLJgdOLFwHUo7L1Dkk4QfsybdRH4ObVxd8509XmKYP
QaYnWRRJc5aYPGyI3LyohpUJdZL+pUGh7Bf9yHbi7AYvqJOW2Q2lxnbtYS3b8+44+GTi5SR7W4wc
il+UulSN/b+xuYnHO1kjpBoL6cVD4///iEl6Um0beKdi8hRbtCUJG2NXnfLFIT8pyhvkP/g4QC8k
08avSV3PRLa4dPmglm0S4NE/wqtyGQ7w4sDOYcyxKfslJ8rUlhReDo1eA7TKgIZvh2+mQaXvSMw+
btj4vAGt76ryRo0sUiiqrung1B+1HBd6iu4flKorfLxdCqGGBQDOlE6JO/+wt4XU43iGM0K8pmwo
nYlzruuIR4XQ7Knym+JIuj+NKQBK+vkTV0+BVMtIuE8yI9T824c3jj3bavZSmNpKrTI52cl8QVI5
vCIfeh3KzLUkIvnovbFlJ1gQUChT03ED+/b25iMMWwGPhUjfyVpte23RRRoy8SefTsapj3s0wfxl
SgrEyKy9G+51vNI7QHnafQ+sHHbYyCUVcIh32jwxqHrwOaj4ilLVSw6uUqVdq4pXwM8qS+y0Qy2S
2XfubqPgW7YgnsttjHHpf9TMkElwReOsNg8uYb4RVAH6oQ+lbpS9i2K4YI9/4dFm5sK+PclAQQ+N
XItfWa/q5/aX9eZ8eMANNs3IW46y2Z1zjmvVwHW7PjOYYuXG3RikT+YVA7eT+w7yY7W3yVU94W09
wemB4Pon8DG6qHhUYAsJR34ExQVgqakmcz8E5uvWZhXQQ1Egy8BtnQJl3UGO1iHxrV17a8u3vC7A
ne2Ep676MuQN/85WH0g71l2okNz1bgZTqXqwz+721yY6G7f2T7USvPHAQBLmri4jzQcwWLwirqdk
teo/sZRF0hhxoDIm2WZe94CTZNj/Rs6Bat7snL31ayZx7S/r4pkRbfkAJ4wgQoAoC4F91RZqEQ3F
FkL3vQmfmarVh/L9X0V2tmICcF245n4CJZYnzeAi3s7LcH1Ug5jk/qJ0j5lmaKfDLwCoy9pvOoQT
piOsBxDrlYZDMdqyRTtnr1UtozJkgaYubix2ton/aZzjJLOlPjWY5Io9T8MJVvek7l39LlDMJbCc
Hf6tgFDicRcpwNQ9KYeHUEE5fPGEey9rAl2Po5UXM+RHk8uvLppp7x1DVLdldznuY5dkh6vUTv9K
mwzsC3wiXgZpIl5oHrOSnIHiBUQlQoWdXojs+8KW1iIpOVVGwCmaYOloBoP9CxN99cbNqyCSg4tS
EAsI0jfYiV/dyN/JN1BAEajUiEL2RKAdCCzBqLiRAsA6BcRpSOtYd1BYifQKZN1afBpnTO2yOfHy
zmNcNqoWsHcY4mhcoeiiU8SUcBCUTg0Ci3zKKz555MfFX4t8Pa/fBXSOOozx2E2jpvbVzckUDGcn
GG0QE9Pl6X3ZfpZzcyhIKh6peOS/9Yw14nzPIon0UGWN7GmDM2y+eRd1tLU3fnkKdxgIQLxP0jcR
wqIG5k9xclWtqPFaORA5OVOm+JEtBK+9zA+Uu6F6rTxV9S5/WkRYzrTzHEys4HUv/iOYaqLIlDou
3RuXymFKbBXXkLF75PRPxCYBUBiFNZSQvSzmMj74boJ192Htx2xMx/L2u4Tpb7s2Du+lgkCs5/Sn
kxXmSonixPhO1OVTzBhN1SmXE8IMZuHg0V0yTrANcc0efc3Pq6vOhgCb1wM97ped13euVzYWLvCE
txXvyMOlg24aQ6lKDrkO+/J+GJeUmdawUOTz0en6L/CoyJhW1389mqOnoKnZx6A02XswPRgiV6J5
b7mhYzTZ378QzLik9MYF4b7BLiqJuZ92EHE4+I9HQbVv5vGV40GkY7PyO7BQDpjhkmBX0BHFbtL5
aeobg4UP3ogDKUm1NFNKazCP6wNv+AChQqgA64T3jPB6hzg9zwnRsiWfeQvmtUa8l7VR6FAlYXvW
p5DeJ1lD/I225iDFenzI+4XJNAuKwDLTZRHo1GF7/iQtHmke83Q+l1cJzTa4CbqA/jkAN8ku5iBG
GTZCFsz7rkW5V5Vt2d+oon5YsJmIw1j2wnKM7myNaB2DOYhArhd6q92Dze0AWfA0wTLRI0ctRMSQ
Ya5X7Dz5aPCEuZ2O6YIgkWr1Kp1P4rfITJiefY+UyAoZPX18VkYzDJtV3Gnhe3wThmf8OkvYL24w
p0WeIrZqNx/X4zXAbOXLt40U7oeuzzdvQ98Yq4iRYLGtanlcvFDEP5hgKALySCL62xFmtr7tSHzF
jeGwPEyFW26ASvgSNZ3G3AZKLf481DQCuo44jZvJ5v6NJE1ufxzYsLxdHofWWP66mw9Xk00p7CYe
qDQ+GeLpWFllEpFCkxbOid4Np5Ky42Z+BGcqQ/OU22Rm1ZAbKtI9C53wxLP3k+y9O/gfCysSGCCT
kCd0a5TF1Djbe7DsBGY05hik9kB34ylhXckBL8QD8paPHFqg7GBAI43uXcTaZhl0d4dtknYlf+s/
xCS4Q/Et5In7geOhYFv8iPywh0cjb+HseHK+ByShM9w2mkJC2BhSJLpIpYLKkvvU8Jwh/Z/TcmT+
MWL6xXt+n7M2t4prAG4STKHlp/VaOUvN7+ku9XkD2bhheUZxCQcshAgVhPrvq5jedV9K341F1F/O
VF/n9+g1oepqtBLP4H6+7tTTpjan7Qd8+1MB05G/RCuMJMK8SqDfOaWFpxiAURWL6YoWLRaIt2K4
mpI0pNNdawgW6413tctbH+b67NGhs76d68xSFWD//IVck9dGpW73AFEX0nLY0LPSuVsnhf8suy+5
/bKvTkb2lW1ctIVsGqU1ylaRDzj0MX1woUyPZB6m+PS/oyaUoRGzeeYFNzKAkb8DUlNn5hk7JjTj
a5vounDFbcyb0qVl+X9Qci9i+XmQ8OBK9UaYUeDGfaUPwlEYZ2vL0nUFxkWNxmV6XZBdpvhdeG9I
CtIWUydGppqOE9w5sjoZT2BoNwYwhek2iIjZG3JHJwytEJ1YpVaub6CaeI+a/hMxKOwvKJGdPg+N
r3CIwphvLZWqZTcCmnlLnNHbwOk8e6+fXY1FKPDnjU/wpIAnwPIrVfASN/RKmTgHQrsxDxAxuIDn
veB9ev5Txmbn48HIivDUJgZ2svoSmguYvqYUDvCR8w00XXJI9XD9gv0HsdB8B27nji1Ns6QkIxnh
TDoeyOxgFT92hY45/K273FMZOYSucf1N7N2KCjrXofMrvZdvHAe2foMoyomsZmdkFnvcameqixXy
WSWQU8J7gh1mZWCeBArXl9FpZHy+0/5wT3opA61updEwYH00sWfLbfzA1kxYI3fqy90PTVMxc8IG
p7ryF6ZzbkyGWlrxL+JGEcCN2CRW2t+NlsUueRr1h2umSG4/Wgrk2fLTqHBr+tfc1qnEngMhVGBl
3uqwLjBSXcqRohNBgFgzXeFXdvD6lXmBdZ1rzectZAEUmW11qxqCqYIgFFTAJIWShBGVLJ1Cd6uF
rsYSy9IbMN3FLL+5vCGviZypGzrBAq2jF916PkWG+//V+9HV5bu/M8k/Xv3ZK3lFYy6qBDVNV/eA
4IgWFO3lXNB/7XIV1TcWFdOeHO27FHO7pNdjNtE2ZL+UyKOlP7089/6bxx+U2udwxZhvsD7raHdQ
BXDEwHbPQJDp3SjnVpgLJz1RqBB0JVOAMVwfoi0yxzOP6NpcFTtdAk2JNQaIxRijopLnGKo4IzuJ
VFROX6F49EMFsdPPzORJdSfG3iuP+fc4HGI2nps98MrB5AX4WqSqOValASgJ0njrmUkqBttH6TDz
p5wVj1kPyb//CrGFA5HNOKAWkASZI63SkVTRFgZvlWzCd1kkHo2bmdkEJAy6DZX9ZVTen0BjlZ66
8CPABT1EUHCUsC0krzCfjYDqCHHThMdqF33/NRUiPA5pzwlLdFXB7x1CeruZpv5jUCBz8+2rr17m
IcjUj2F4jT//E9eUnO3Xb8MVbjHPsH6zk7AGNw5rqpBjCj7inbEJqCdx6Qg3yEPNLUdpUK63pplL
Tv5AHQmqHt8m8vSX7o481PsAoY2gpOR/gCf+Ixj2oGQT9G4vY7DHDfmC3ULx6XNos4jM9bLaAZn9
mziD/1mPLnOPpi8ree6RYxZ7IHt99KmviUy9m2PG0Sm8fuT9nPnJFWdLDoKIpOm6w1pw7hGYZE7W
5cMt4lUtAQQzgTV15L/6BkeycrEIsSLN8knsusk+g5GgQ8+CHsQJsdc00Hre0DAcitwSfLiUv903
Y+r9Tjb4EK6Jws1+xt4jpxISpHewBhmM7qJ5C7nvj7FCmdsBwp/ApciRwaji5D6OiNVYABlTkDWM
8zePYO/ww9UqCTvx9QQvveXYGhxc/1hmsvOhKS2g8GHwPoCgviPK65Dk2G+/Aqh/+k/QopdvrHb0
SDQkrZFZ7kDMVXxvafNJVK1jB1DOIuAHfAVnzSL4jUoB8XBsP3CNMFpsHBdhkZRWoZ8MyO2KIDHZ
JXvGPwPRzZVrQdqXTjycRNXglk1qkHR+XvxTiBypkqN4eP9oz98if/q+vkLgKlA2+vL+Jmer+EzP
/6abbvihrFitsWN7NLBKwl4H23F12nj+2Ah1rBdkEP6L4fr61Wt7ubf6gw6XARJpk5KsblboklM6
aYLWeyLeTFjq9i8OOemv2soWT6pUG84z6T0CL/PzCN2/1A9DrBpPz7eNYvQmkyjb31lZ+sWdtJy/
2esIpsFwktRNUwUojbCwV0Tv3kWSefsPJ9sLZAIzahnBUcOVmxEhtBSjTS3V8NcDANdHOsocFGNA
XW7AESvtXZieqvjMPLvtos8SO0FCQ+A0+YX2hgzu7eCq4AznXhIl39b3V8Axq1fD6x3CQQuYST0w
hC6cAcgGo25g8IOXkfUKGXujuLOy+Uzr4XNtwmQ2QO03bbXC7VE9+TbsxlOt5kymMKZBLEXGLYwl
cOtOR93KHF2rwZ9ellDHNUHBrM2Ltjrbub/5/O7671q8pNMZujF/r8s8Z2mz7GTxcWX+GGDO0Lq6
SHLIbqbRRkU7uaG8LrdhOdLUHbyTdITlegC/fsTEG6iyQUZ2hv143i+d85ZlrzcF2KYZA8Twb3On
FanG8rLpwHUf34ZSJa38eQ1+yZ9w+pejQVKw6wz405yCIP9zLmX/O5gppOZInBKG3R5+21GSDIHt
LnQb1C2w7bbRLdbkCCzU7MHh5b9aez2dCDlz1NPer21VOSwSQlvxtepH6LDkiNvn64r9sP3FSKHq
3Z0x7YKe/+xsotO8JnQ4HKxuk2GuNTH/gIv9CVCCEqIKGET2VGXKz5NI4v/kCO4c6zSwiGYUG4gZ
tDmLUHBvxFKenR9OyhqNHaMsOTRm0XOim6PpghWsp49jGFXfb4LNqXHa+Ytyzzx+ftL4BK85cXgl
RFYx6qNdoWOcAUEWvzRHpkxqcv25hsLT+QqlHel1xjV9cGoAFTic946jo16Iks9scuqJrrxs0j3w
SiJ8gcmNQTat+W2DQ9i5s2aLhC0Hf/o2w9P5WTMhGAzDrp/nPqRIDCc102m+IApyyimIz3KSKIBS
aFHSp761XRKI3bkvXxLhcZKgIJcQF6+7DEPyGCZJiYVLhQpEkYijKNuHC2cdox9A+MW+/zq3xZxs
ZsGMWfU3O6oUumzdcr7MLI1fKD3W3Aj5/JyJ5aGa5zfPvJLgJ1h5QUq7166H4hyxexkDik/36RBt
04B4qeuuA9GviPMmsHzDgoJUDtc0pLoQIAfTTwrjKcPXOmPjSIUOtHm1maXK4rokvyMrVV5Mf2CK
7gmNRnSLEqgClDorRMkAj/Tq16cJulJJI9PV9yc5lTqK2IuOn1edxsZKPHScT784tbX2e3tVAOIO
ZKxPUxOvu/bbA6B8vQ8VkzJ6u55C/5ggp8/bRbBn89To8jKQ0SfX7e0OMqFCpXiNrXsR/N8P/Rva
5f9D5ybQ49qBIl7f7X0NKtQNo/WilFg58he1EuIFRsfvz2CJSAPyzqFWGDuW46zw3HTpp4mdcAIN
wFhxb9VjgvnbzLyF0tKh8IvrmfU6sDzLFWboK8fLrKjuiZOED+C2AB32zBMYbdgangIxx+uJBHN8
sKvY6LjBYVapCJ8ujMd3Xi151ORWJRQkU3u53BhBxWsaGLOTl0TCnYxi5rcpkbynNm07Nb3rBPQx
iUO0Qpj6ovfvil9SxrfSHvGs5M7kGXQk57Jc02jyhOq8zqSpsUnjEVj1r4Hr3mcuCCTMJwuAmTSf
gMEi+tNU4LP4FTM/LFn4U/qOz5saOhYm6mQCXJs3yEzulu86ptOK9y8PNngKZQAokuwrRZAZDzXp
g76ukoW6qgqCWeIm6IW9L/44wzPiL4GP91zqEKXnad3A1bLK8DPoho71pDcHdH/DIJW4R3kegbbA
2CNeWNuyCLyFWuTuseAWft0+X2orplsp7j2kxRQi1q1Q2QumWvYqm55OwE60LXv3bAaL2Fp2Ji4u
Iz3ix//QUlOAHPE4DdLupftVsmRpaZ6uoNegvM5YajDnwecLL1kf6ZrzwbpmiEMXuqV48Qgtzikw
ECDABiFmBXp7hon6EcxNGTtL7QemV6tOscRgFaj7TU2hn9z2Qa5sf0rUrx+70dgHv6/6AW2ZPCpn
tLdLAejRQNOeGW/gSjo0HkA6HGiqsAaeeGm37rIF150s4RoH4+ayyAAvMVys9ApuRjLUVuICYJp/
kBoc088fMadMZyIHl4DY50CerVtjOxB+0d4+w3/A8xL4oRKJE2u503t8pMMoxJMxzpuu0IqQ5aVO
SQJLNlpDmw0mf0UYK7Z6PUbSC81FtwQjxb8cmJnvp4dRWWVSailw+3n+aIzBEOIJq8+zq5iVXs+c
5kiLVz0CEXAIuyoNt1dpEidIm91nSozkJ81/xJ1riIBGefgj64Y1owu2r4snJosk9BgIzUwrwxkK
OXVRl2wSxuI+ueaSBO+9LrcFv0ibPQngYxkGtc55AhZZ3jqJxNIhLG60lgAkcGJPR0gRL0zgH83Z
SMZR+ZOrOlGZDhOtwKYqCvtx8ExqRUY3Q8dBY7w7eZU5ur/VskbL12CRj5CD9GRkOq5VfbBkUamC
kKsVza7u14jTZrLCPaC5gZPRot/ithN+fMlAPWjNqxeTC6WqIOtVWkInCOJFAtdXeTuTNi9eZqSl
WSAfoO7G4sRRCL5cTavONRhTSDLNEEw6puw5DAbxhrdlWnEj+N8KbUBw9+in9/STg1n6pppXoRR/
1S6RTntKugGGW/G1G29D5MZnGADkDx5TVO3o4R/2DqLBUForpf7AKwbYYAgmzg9GMjA7QqCPOw+g
YTzzTo22I7X6pCVoWj3ECOP+iqawQjD+bvsUQ4+uNuaJynQ+XeMAiD9sbdpMOOJT5OAvGcvsbojy
ygco7bp5I+B6KGTDiJgvq2UCAbl+QlNfa+d6I5AngmMVMB1smKyESot0ib1N4lOXZF5KMCfk9LbV
UCOT7OsDFWQKwVNpcxV4ga8yrIJcN6IJQCXs5ZYadu7TCPdelSqYV/9RfLiZWZZcAf4LS01jkB19
bj77GLaeDFUm72CnX3/CzMwVT0hpH//4bHm0MOfePuNeoV1wD7W6ExQCoyvxtO10p/rrW0vOPT7z
+kjN7/g9h9LE+FLXh36JbpfBFWQlIv6mbA+izlXoXGrM7U+GvYZipqA8IX4jPUgmiIrpzd9i6QZu
2Zh5JAolwqr/xI5fnsMT5Gw5GZiVQUNMU/2gew+fQHL3x9DUlCTpJ/upaegKChHc8ipCBBHx8jrO
86G3DNdnxHYLmjCATNNzyzV+uQbDjT2cnzCRIRpmrjPEckqrb0pJFyzFOP1eIhy+1eBTNJfrqfIi
xmic40CU6rda9mj20TIRHr5JRSn7cPBE5lNlm+TwlNYAKkSIXGZxvNlaVFyUm9VKHQ5HMIC0SNaW
znelTs2roO36QsdOea50hDRWqh920AzGRn9uhQ1ghZmHhMD+KrS/TGMwSrvnEe0zcDSQphHowck8
0eH1xGNKPuSfGxj/yLjM0c3/hNxEDbM9JqIr+Wg2vTRo3ojPLT+UKXyiO3yqrOj3QNiuY+kd4Qou
lmzldTt5ClslyCyAoCtb2Zo8nFKWGmiRGJTnkD3HAo7V5U9EsJh2QlSzIzc9VyBGIADO9K7sIqLV
Et4TXzrqvaavEl89aWj7FG2UmZcPfD9Zb6bHsBhh2n16NayKZlU12Jn9JlLI9NED8OPRaTYw1V/y
qL1Af82B8Kri8OC/rf44ceMb3bmkRtyYx/8zTW8udKSFt0Uhh2tZSpHv9VvFgq6v3V/OAgSwHwlP
yGSr7m4FqsRt6wyKKoFeBPtKidPX764PdDAd0VE95PNhpKApT9x4KwDddq6OCTNXW8ssKfq4AMvM
I8I8x0oFXoZYLoRPzAWM63TICNCl8PYQeUg8BadeWA3W6vNKOuHmz9me9gu1qWvB/B4yWjB4Zw85
0QOMBGYdi4u/lUbGnkARnJWYX/pjW5fEv94CRopbjPYxl+GRwJECsX9ItYPja9lg/Y/HPDlVwrVj
gEYhwih1unHxnPa3WB+C8i/Cfs+ho0wn9yNKBT3zuXAj5nJgjchfbT2OdouRMpGbkosTh+q4Bibl
inp/BugIX0QExdw4lrmY4sAiT+/hEHUAVUVu+U8yibGPhfQKFF660vbBJAHQqFqS2sOzmJ8v3FBS
90AUi+2A8Eg4BdgfbTaeFKXwDsmF6fw+xwqpGERPvIXq2scVv9G26CS0ZvDAwoo9m+YdmtxXKrLk
PXWfjzX2gSyNsV5s7Di9mQYTWo9wH8o9RDoVEuoaKvt1kV5RAvc25gD5EnCgvRLo3iitdsWwB+BD
ZuNF30BYJS34bVLhEWVMyG7GkIq49mK2ePULzCMpzKvrPi81o0A4woW5YrKFYTvRp0CDVQ/GRC2V
qKeVeDlnku7ScZhgxc3Fw8ygZZAqi605RKNJAXrjctN8/s+Xo6LAM+arRa8AR+8waOW4+wbf5NmL
RammQfAmyogMEoeYFjnABVkAXO94N5kbMSIPpBODa/ZJPXrEUNYrL5RYcakhgCgXymWq1KFE9awC
UR0R6ueRRzNTTYbvfrADSGY4kZnwklSqUg0a+CI43hwjgGgFuRKKUjm9o5PvSh3VPt9K9eClGZ82
8cU9xWje1B2BorbjjJ1yP9eD/a8ue6bA5NYEoA5+DGhHy/Y7KXcnV0r0FgvB/9xxzA8z2r81ydEG
/f5iE1pdTFAUyYG1ojKGdpPSwARMxH5S1pZo/d5esrDZUrg9ZmyrO/gu94RaLbUgaK16CiD7A1TY
aIWgO3fkmAtx5IUNLKo4Nb9c84mchKF3TPnkpLI4VUDsRvfOhpEGNNoWpg0D3UK315uTNNLSu9TA
0HsR9zGtn7oZz8KyyeR/TDZKnUUdpYa8L0Zts7tWdPWLWaq3w4iBZjL7CmB0dTdhTbHLqsNm8e6E
Z8I0FcTq6+InXE6+0SIUOGwWIBz3i3wH5je0uHTZfQx/MP+6rdQVw8MmMTydagtUNGDhn1Nl9JU4
weBl3ElcigOujGr3lKSl2rpRNNVAFEfDSew2kAURguOtKVJw7E6fvo7R9mfLQ2wd41zBZexdUnf9
TYU1iC7O0rIAoHoh5/LVpymGkYaJdhDgrUJZLDAqK5DXBE1ANDje/bc1HifxOCb4Jhr8AO+h/c1l
Lzk0KLe5eZwLpW/NpYF2PJKYFNIVombZ5l6VJ+Rfnd5xNux04EGMq0FRtkNP8QMiIvUfqU4uvp8h
hiI1ZrCNdpFjhSLSkjQVQeq400tQ6nrf5b3F8rGJpnJtytmH6wmNN28eDa+oSDUvjtNYJjNoJ0+c
fFiPLygUzpe8Oup1VFGWkdaUh3eCO/unFff8Tu/4qoHJU2XYiswF7XAHQMihnPLIto5qFUhgFpJY
vOp4VNxasB210FgHZNF1jWFMI6vu1qTmNGsndHQR5twVUS2+lQP+I1n3YijEWtQ3hqO9Zom56fWy
jlRzRQafwl7Pb1fH+HeoZnIJGXdf
`protect end_protected
